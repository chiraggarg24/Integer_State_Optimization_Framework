//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-10-29 20:45:32.425445
// Design Name: vanilla
// Module Name: sigmoidLUT_in6b3p_out16b15p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 6 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in6b3p_out16b15p #(
    parameter PRECISION_INPUT_BITS = 6,
    parameter PRECISION_OUTPUT_BITS = 16
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			6'b000000: sigmoid_out <= 16'b0100000000000000;    //sigmoid(0.000000) ≈ 0.500000
			6'b000001: sigmoid_out <= 16'b0100001111111111;    //sigmoid(0.125000) ≈ 0.531219
			6'b000010: sigmoid_out <= 16'b0100011111110101;    //sigmoid(0.250000) ≈ 0.562164
			6'b000011: sigmoid_out <= 16'b0100101111011100;    //sigmoid(0.375000) ≈ 0.592651
			6'b000100: sigmoid_out <= 16'b0100111110101101;    //sigmoid(0.500000) ≈ 0.622467
			6'b000101: sigmoid_out <= 16'b0101001101100000;    //sigmoid(0.625000) ≈ 0.651367
			6'b000110: sigmoid_out <= 16'b0101011011101111;    //sigmoid(0.750000) ≈ 0.679169
			6'b000111: sigmoid_out <= 16'b0101101001010111;    //sigmoid(0.875000) ≈ 0.705780
			6'b001000: sigmoid_out <= 16'b0101110110010011;    //sigmoid(1.000000) ≈ 0.731049
			6'b001001: sigmoid_out <= 16'b0110000010100001;    //sigmoid(1.125000) ≈ 0.754913
			6'b001010: sigmoid_out <= 16'b0110001101111111;    //sigmoid(1.250000) ≈ 0.777313
			6'b001011: sigmoid_out <= 16'b0110011000101011;    //sigmoid(1.375000) ≈ 0.798187
			6'b001100: sigmoid_out <= 16'b0110100010100110;    //sigmoid(1.500000) ≈ 0.817566
			6'b001101: sigmoid_out <= 16'b0110101011110001;    //sigmoid(1.625000) ≈ 0.835480
			6'b001110: sigmoid_out <= 16'b0110110100001101;    //sigmoid(1.750000) ≈ 0.851959
			6'b001111: sigmoid_out <= 16'b0110111011111011;    //sigmoid(1.875000) ≈ 0.867035
			6'b010000: sigmoid_out <= 16'b0111000010111110;    //sigmoid(2.000000) ≈ 0.880798
			6'b010001: sigmoid_out <= 16'b0111001001011000;    //sigmoid(2.125000) ≈ 0.893311
			6'b010010: sigmoid_out <= 16'b0111001111001100;    //sigmoid(2.250000) ≈ 0.904663
			6'b010011: sigmoid_out <= 16'b0111010100011011;    //sigmoid(2.375000) ≈ 0.914886
			6'b010100: sigmoid_out <= 16'b0111011001001010;    //sigmoid(2.500000) ≈ 0.924133
			6'b010101: sigmoid_out <= 16'b0111011101011011;    //sigmoid(2.625000) ≈ 0.932465
			6'b010110: sigmoid_out <= 16'b0111100001001111;    //sigmoid(2.750000) ≈ 0.939911
			6'b010111: sigmoid_out <= 16'b0111100100101010;    //sigmoid(2.875000) ≈ 0.946594
			6'b011000: sigmoid_out <= 16'b0111100111101110;    //sigmoid(3.000000) ≈ 0.952576
			6'b011001: sigmoid_out <= 16'b0111101010011101;    //sigmoid(3.125000) ≈ 0.957916
			6'b011010: sigmoid_out <= 16'b0111101100111001;    //sigmoid(3.250000) ≈ 0.962677
			6'b011011: sigmoid_out <= 16'b0111101111000100;    //sigmoid(3.375000) ≈ 0.966919
			6'b011100: sigmoid_out <= 16'b0111110000111111;    //sigmoid(3.500000) ≈ 0.970673
			6'b011101: sigmoid_out <= 16'b0111110010101101;    //sigmoid(3.625000) ≈ 0.974030
			6'b011110: sigmoid_out <= 16'b0111110100001111;    //sigmoid(3.750000) ≈ 0.977020
			6'b011111: sigmoid_out <= 16'b0111110101100110;    //sigmoid(3.875000) ≈ 0.979675
			6'b100000: sigmoid_out <= 16'b0111110110110011;    //sigmoid(4.000000) ≈ 0.982025
			6'b100001: sigmoid_out <= 16'b0111110111110111;    //sigmoid(4.125000) ≈ 0.984100
			6'b100010: sigmoid_out <= 16'b0111111000110011;    //sigmoid(4.250000) ≈ 0.985931
			6'b100011: sigmoid_out <= 16'b0111111001101001;    //sigmoid(4.375000) ≈ 0.987579
			6'b100100: sigmoid_out <= 16'b0111111010011000;    //sigmoid(4.500000) ≈ 0.989014
			6'b100101: sigmoid_out <= 16'b0111111011000010;    //sigmoid(4.625000) ≈ 0.990295
			6'b100110: sigmoid_out <= 16'b0111111011100111;    //sigmoid(4.750000) ≈ 0.991425
			6'b100111: sigmoid_out <= 16'b0111111100001000;    //sigmoid(4.875000) ≈ 0.992432
			6'b101000: sigmoid_out <= 16'b0111111100100101;    //sigmoid(5.000000) ≈ 0.993317
			6'b101001: sigmoid_out <= 16'b0111111100111110;    //sigmoid(5.125000) ≈ 0.994080
			6'b101010: sigmoid_out <= 16'b0111111101010101;    //sigmoid(5.250000) ≈ 0.994781
			6'b101011: sigmoid_out <= 16'b0111111101101001;    //sigmoid(5.375000) ≈ 0.995392
			6'b101100: sigmoid_out <= 16'b0111111101111011;    //sigmoid(5.500000) ≈ 0.995941
			6'b101101: sigmoid_out <= 16'b0111111110001010;    //sigmoid(5.625000) ≈ 0.996399
			6'b101110: sigmoid_out <= 16'b0111111110011000;    //sigmoid(5.750000) ≈ 0.996826
			6'b101111: sigmoid_out <= 16'b0111111110100100;    //sigmoid(5.875000) ≈ 0.997192
			6'b110000: sigmoid_out <= 16'b0111111110101111;    //sigmoid(6.000000) ≈ 0.997528
			6'b110001: sigmoid_out <= 16'b0111111110111000;    //sigmoid(6.125000) ≈ 0.997803
			6'b110010: sigmoid_out <= 16'b0111111111000001;    //sigmoid(6.250000) ≈ 0.998077
			6'b110011: sigmoid_out <= 16'b0111111111001000;    //sigmoid(6.375000) ≈ 0.998291
			6'b110100: sigmoid_out <= 16'b0111111111001111;    //sigmoid(6.500000) ≈ 0.998505
			6'b110101: sigmoid_out <= 16'b0111111111010101;    //sigmoid(6.625000) ≈ 0.998688
			6'b110110: sigmoid_out <= 16'b0111111111011010;    //sigmoid(6.750000) ≈ 0.998840
			6'b110111: sigmoid_out <= 16'b0111111111011110;    //sigmoid(6.875000) ≈ 0.998962
			6'b111000: sigmoid_out <= 16'b0111111111100010;    //sigmoid(7.000000) ≈ 0.999084
			6'b111001: sigmoid_out <= 16'b0111111111100110;    //sigmoid(7.125000) ≈ 0.999207
			6'b111010: sigmoid_out <= 16'b0111111111101001;    //sigmoid(7.250000) ≈ 0.999298
			6'b111011: sigmoid_out <= 16'b0111111111101011;    //sigmoid(7.375000) ≈ 0.999359
			6'b111100: sigmoid_out <= 16'b0111111111101110;    //sigmoid(7.500000) ≈ 0.999451
			6'b111101: sigmoid_out <= 16'b0111111111110000;    //sigmoid(7.625000) ≈ 0.999512
			6'b111110: sigmoid_out <= 16'b0111111111110010;    //sigmoid(7.750000) ≈ 0.999573
			6'b111111: sigmoid_out <= 16'b0111111111110100;    //sigmoid(7.875000) ≈ 0.999634

        endcase
    end
endmodule