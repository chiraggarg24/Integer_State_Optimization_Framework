//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
// 
// Create Date: 2019-06-28 11:46:00.454444
// Design Name: vanilla
// Module Name: sigmoidLUT_7bit_7point
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 7 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
// 
// Additional Comments: Generated by LUT_generator_sigmoid.py
// 
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_7bit_7point #(
    parameter PRECISION_BITS = 7
)(
    input[PRECISION_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			7'b0000000: sigmoid_out <= 7'b1000000;    //sigmoid(0.000000) ≈ 0.500000
			7'b0000001: sigmoid_out <= 7'b1000000;    //sigmoid(0.007812) ≈ 0.500000
			7'b0000010: sigmoid_out <= 7'b1000000;    //sigmoid(0.015625) ≈ 0.500000
			7'b0000011: sigmoid_out <= 7'b1000001;    //sigmoid(0.023438) ≈ 0.507812
			7'b0000100: sigmoid_out <= 7'b1000001;    //sigmoid(0.031250) ≈ 0.507812
			7'b0000101: sigmoid_out <= 7'b1000001;    //sigmoid(0.039062) ≈ 0.507812
			7'b0000110: sigmoid_out <= 7'b1000001;    //sigmoid(0.046875) ≈ 0.507812
			7'b0000111: sigmoid_out <= 7'b1000010;    //sigmoid(0.054688) ≈ 0.515625
			7'b0001000: sigmoid_out <= 7'b1000010;    //sigmoid(0.062500) ≈ 0.515625
			7'b0001001: sigmoid_out <= 7'b1000010;    //sigmoid(0.070312) ≈ 0.515625
			7'b0001010: sigmoid_out <= 7'b1000010;    //sigmoid(0.078125) ≈ 0.515625
			7'b0001011: sigmoid_out <= 7'b1000011;    //sigmoid(0.085938) ≈ 0.523438
			7'b0001100: sigmoid_out <= 7'b1000011;    //sigmoid(0.093750) ≈ 0.523438
			7'b0001101: sigmoid_out <= 7'b1000011;    //sigmoid(0.101562) ≈ 0.523438
			7'b0001110: sigmoid_out <= 7'b1000011;    //sigmoid(0.109375) ≈ 0.523438
			7'b0001111: sigmoid_out <= 7'b1000100;    //sigmoid(0.117188) ≈ 0.531250
			7'b0010000: sigmoid_out <= 7'b1000100;    //sigmoid(0.125000) ≈ 0.531250
			7'b0010001: sigmoid_out <= 7'b1000100;    //sigmoid(0.132812) ≈ 0.531250
			7'b0010010: sigmoid_out <= 7'b1000100;    //sigmoid(0.140625) ≈ 0.531250
			7'b0010011: sigmoid_out <= 7'b1000101;    //sigmoid(0.148438) ≈ 0.539062
			7'b0010100: sigmoid_out <= 7'b1000101;    //sigmoid(0.156250) ≈ 0.539062
			7'b0010101: sigmoid_out <= 7'b1000101;    //sigmoid(0.164062) ≈ 0.539062
			7'b0010110: sigmoid_out <= 7'b1000101;    //sigmoid(0.171875) ≈ 0.539062
			7'b0010111: sigmoid_out <= 7'b1000110;    //sigmoid(0.179688) ≈ 0.546875
			7'b0011000: sigmoid_out <= 7'b1000110;    //sigmoid(0.187500) ≈ 0.546875
			7'b0011001: sigmoid_out <= 7'b1000110;    //sigmoid(0.195312) ≈ 0.546875
			7'b0011010: sigmoid_out <= 7'b1000110;    //sigmoid(0.203125) ≈ 0.546875
			7'b0011011: sigmoid_out <= 7'b1000111;    //sigmoid(0.210938) ≈ 0.554688
			7'b0011100: sigmoid_out <= 7'b1000111;    //sigmoid(0.218750) ≈ 0.554688
			7'b0011101: sigmoid_out <= 7'b1000111;    //sigmoid(0.226562) ≈ 0.554688
			7'b0011110: sigmoid_out <= 7'b1000111;    //sigmoid(0.234375) ≈ 0.554688
			7'b0011111: sigmoid_out <= 7'b1001000;    //sigmoid(0.242188) ≈ 0.562500
			7'b0100000: sigmoid_out <= 7'b1001000;    //sigmoid(0.250000) ≈ 0.562500
			7'b0100001: sigmoid_out <= 7'b1001000;    //sigmoid(0.257812) ≈ 0.562500
			7'b0100010: sigmoid_out <= 7'b1001000;    //sigmoid(0.265625) ≈ 0.562500
			7'b0100011: sigmoid_out <= 7'b1001001;    //sigmoid(0.273438) ≈ 0.570312
			7'b0100100: sigmoid_out <= 7'b1001001;    //sigmoid(0.281250) ≈ 0.570312
			7'b0100101: sigmoid_out <= 7'b1001001;    //sigmoid(0.289062) ≈ 0.570312
			7'b0100110: sigmoid_out <= 7'b1001001;    //sigmoid(0.296875) ≈ 0.570312
			7'b0100111: sigmoid_out <= 7'b1001010;    //sigmoid(0.304688) ≈ 0.578125
			7'b0101000: sigmoid_out <= 7'b1001010;    //sigmoid(0.312500) ≈ 0.578125
			7'b0101001: sigmoid_out <= 7'b1001010;    //sigmoid(0.320312) ≈ 0.578125
			7'b0101010: sigmoid_out <= 7'b1001010;    //sigmoid(0.328125) ≈ 0.578125
			7'b0101011: sigmoid_out <= 7'b1001011;    //sigmoid(0.335938) ≈ 0.585938
			7'b0101100: sigmoid_out <= 7'b1001011;    //sigmoid(0.343750) ≈ 0.585938
			7'b0101101: sigmoid_out <= 7'b1001011;    //sigmoid(0.351562) ≈ 0.585938
			7'b0101110: sigmoid_out <= 7'b1001011;    //sigmoid(0.359375) ≈ 0.585938
			7'b0101111: sigmoid_out <= 7'b1001100;    //sigmoid(0.367188) ≈ 0.593750
			7'b0110000: sigmoid_out <= 7'b1001100;    //sigmoid(0.375000) ≈ 0.593750
			7'b0110001: sigmoid_out <= 7'b1001100;    //sigmoid(0.382812) ≈ 0.593750
			7'b0110010: sigmoid_out <= 7'b1001100;    //sigmoid(0.390625) ≈ 0.593750
			7'b0110011: sigmoid_out <= 7'b1001101;    //sigmoid(0.398438) ≈ 0.601562
			7'b0110100: sigmoid_out <= 7'b1001101;    //sigmoid(0.406250) ≈ 0.601562
			7'b0110101: sigmoid_out <= 7'b1001101;    //sigmoid(0.414062) ≈ 0.601562
			7'b0110110: sigmoid_out <= 7'b1001101;    //sigmoid(0.421875) ≈ 0.601562
			7'b0110111: sigmoid_out <= 7'b1001110;    //sigmoid(0.429688) ≈ 0.609375
			7'b0111000: sigmoid_out <= 7'b1001110;    //sigmoid(0.437500) ≈ 0.609375
			7'b0111001: sigmoid_out <= 7'b1001110;    //sigmoid(0.445312) ≈ 0.609375
			7'b0111010: sigmoid_out <= 7'b1001110;    //sigmoid(0.453125) ≈ 0.609375
			7'b0111011: sigmoid_out <= 7'b1001110;    //sigmoid(0.460938) ≈ 0.609375
			7'b0111100: sigmoid_out <= 7'b1001111;    //sigmoid(0.468750) ≈ 0.617188
			7'b0111101: sigmoid_out <= 7'b1001111;    //sigmoid(0.476562) ≈ 0.617188
			7'b0111110: sigmoid_out <= 7'b1001111;    //sigmoid(0.484375) ≈ 0.617188
			7'b0111111: sigmoid_out <= 7'b1001111;    //sigmoid(0.492188) ≈ 0.617188
			7'b1000000: sigmoid_out <= 7'b1010000;    //sigmoid(0.500000) ≈ 0.625000
			7'b1000001: sigmoid_out <= 7'b1010000;    //sigmoid(0.507812) ≈ 0.625000
			7'b1000010: sigmoid_out <= 7'b1010000;    //sigmoid(0.515625) ≈ 0.625000
			7'b1000011: sigmoid_out <= 7'b1010000;    //sigmoid(0.523438) ≈ 0.625000
			7'b1000100: sigmoid_out <= 7'b1010001;    //sigmoid(0.531250) ≈ 0.632812
			7'b1000101: sigmoid_out <= 7'b1010001;    //sigmoid(0.539062) ≈ 0.632812
			7'b1000110: sigmoid_out <= 7'b1010001;    //sigmoid(0.546875) ≈ 0.632812
			7'b1000111: sigmoid_out <= 7'b1010001;    //sigmoid(0.554688) ≈ 0.632812
			7'b1001000: sigmoid_out <= 7'b1010010;    //sigmoid(0.562500) ≈ 0.640625
			7'b1001001: sigmoid_out <= 7'b1010010;    //sigmoid(0.570312) ≈ 0.640625
			7'b1001010: sigmoid_out <= 7'b1010010;    //sigmoid(0.578125) ≈ 0.640625
			7'b1001011: sigmoid_out <= 7'b1010010;    //sigmoid(0.585938) ≈ 0.640625
			7'b1001100: sigmoid_out <= 7'b1010010;    //sigmoid(0.593750) ≈ 0.640625
			7'b1001101: sigmoid_out <= 7'b1010011;    //sigmoid(0.601562) ≈ 0.648438
			7'b1001110: sigmoid_out <= 7'b1010011;    //sigmoid(0.609375) ≈ 0.648438
			7'b1001111: sigmoid_out <= 7'b1010011;    //sigmoid(0.617188) ≈ 0.648438
			7'b1010000: sigmoid_out <= 7'b1010011;    //sigmoid(0.625000) ≈ 0.648438
			7'b1010001: sigmoid_out <= 7'b1010100;    //sigmoid(0.632812) ≈ 0.656250
			7'b1010010: sigmoid_out <= 7'b1010100;    //sigmoid(0.640625) ≈ 0.656250
			7'b1010011: sigmoid_out <= 7'b1010100;    //sigmoid(0.648438) ≈ 0.656250
			7'b1010100: sigmoid_out <= 7'b1010100;    //sigmoid(0.656250) ≈ 0.656250
			7'b1010101: sigmoid_out <= 7'b1010101;    //sigmoid(0.664062) ≈ 0.664062
			7'b1010110: sigmoid_out <= 7'b1010101;    //sigmoid(0.671875) ≈ 0.664062
			7'b1010111: sigmoid_out <= 7'b1010101;    //sigmoid(0.679688) ≈ 0.664062
			7'b1011000: sigmoid_out <= 7'b1010101;    //sigmoid(0.687500) ≈ 0.664062
			7'b1011001: sigmoid_out <= 7'b1010101;    //sigmoid(0.695312) ≈ 0.664062
			7'b1011010: sigmoid_out <= 7'b1010110;    //sigmoid(0.703125) ≈ 0.671875
			7'b1011011: sigmoid_out <= 7'b1010110;    //sigmoid(0.710938) ≈ 0.671875
			7'b1011100: sigmoid_out <= 7'b1010110;    //sigmoid(0.718750) ≈ 0.671875
			7'b1011101: sigmoid_out <= 7'b1010110;    //sigmoid(0.726562) ≈ 0.671875
			7'b1011110: sigmoid_out <= 7'b1010110;    //sigmoid(0.734375) ≈ 0.671875
			7'b1011111: sigmoid_out <= 7'b1010111;    //sigmoid(0.742188) ≈ 0.679688
			7'b1100000: sigmoid_out <= 7'b1010111;    //sigmoid(0.750000) ≈ 0.679688
			7'b1100001: sigmoid_out <= 7'b1010111;    //sigmoid(0.757812) ≈ 0.679688
			7'b1100010: sigmoid_out <= 7'b1010111;    //sigmoid(0.765625) ≈ 0.679688
			7'b1100011: sigmoid_out <= 7'b1011000;    //sigmoid(0.773438) ≈ 0.687500
			7'b1100100: sigmoid_out <= 7'b1011000;    //sigmoid(0.781250) ≈ 0.687500
			7'b1100101: sigmoid_out <= 7'b1011000;    //sigmoid(0.789062) ≈ 0.687500
			7'b1100110: sigmoid_out <= 7'b1011000;    //sigmoid(0.796875) ≈ 0.687500
			7'b1100111: sigmoid_out <= 7'b1011000;    //sigmoid(0.804688) ≈ 0.687500
			7'b1101000: sigmoid_out <= 7'b1011001;    //sigmoid(0.812500) ≈ 0.695312
			7'b1101001: sigmoid_out <= 7'b1011001;    //sigmoid(0.820312) ≈ 0.695312
			7'b1101010: sigmoid_out <= 7'b1011001;    //sigmoid(0.828125) ≈ 0.695312
			7'b1101011: sigmoid_out <= 7'b1011001;    //sigmoid(0.835938) ≈ 0.695312
			7'b1101100: sigmoid_out <= 7'b1011010;    //sigmoid(0.843750) ≈ 0.703125
			7'b1101101: sigmoid_out <= 7'b1011010;    //sigmoid(0.851562) ≈ 0.703125
			7'b1101110: sigmoid_out <= 7'b1011010;    //sigmoid(0.859375) ≈ 0.703125
			7'b1101111: sigmoid_out <= 7'b1011010;    //sigmoid(0.867188) ≈ 0.703125
			7'b1110000: sigmoid_out <= 7'b1011010;    //sigmoid(0.875000) ≈ 0.703125
			7'b1110001: sigmoid_out <= 7'b1011011;    //sigmoid(0.882812) ≈ 0.710938
			7'b1110010: sigmoid_out <= 7'b1011011;    //sigmoid(0.890625) ≈ 0.710938
			7'b1110011: sigmoid_out <= 7'b1011011;    //sigmoid(0.898438) ≈ 0.710938
			7'b1110100: sigmoid_out <= 7'b1011011;    //sigmoid(0.906250) ≈ 0.710938
			7'b1110101: sigmoid_out <= 7'b1011011;    //sigmoid(0.914062) ≈ 0.710938
			7'b1110110: sigmoid_out <= 7'b1011100;    //sigmoid(0.921875) ≈ 0.718750
			7'b1110111: sigmoid_out <= 7'b1011100;    //sigmoid(0.929688) ≈ 0.718750
			7'b1111000: sigmoid_out <= 7'b1011100;    //sigmoid(0.937500) ≈ 0.718750
			7'b1111001: sigmoid_out <= 7'b1011100;    //sigmoid(0.945312) ≈ 0.718750
			7'b1111010: sigmoid_out <= 7'b1011100;    //sigmoid(0.953125) ≈ 0.718750
			7'b1111011: sigmoid_out <= 7'b1011101;    //sigmoid(0.960938) ≈ 0.726562
			7'b1111100: sigmoid_out <= 7'b1011101;    //sigmoid(0.968750) ≈ 0.726562
			7'b1111101: sigmoid_out <= 7'b1011101;    //sigmoid(0.976562) ≈ 0.726562
			7'b1111110: sigmoid_out <= 7'b1011101;    //sigmoid(0.984375) ≈ 0.726562
			7'b1111111: sigmoid_out <= 7'b1011101;    //sigmoid(0.992188) ≈ 0.726562

        endcase
    end
endmodule