//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2020-04-24 09:11:58.477876
// Design Name: vanilla
// Module Name: sigmoidLUT_in6b1p_out16b15p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 6 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in6b1p_out16b15p #(
    parameter PRECISION_INPUT_BITS = 6,
    parameter PRECISION_OUTPUT_BITS = 16
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			6'b000000: sigmoid_out <= 16'b0100000000000000;    //sigmoid(0.000000) ≈ 0.500000
			6'b000001: sigmoid_out <= 16'b0100111110101101;    //sigmoid(0.500000) ≈ 0.622467
			6'b000010: sigmoid_out <= 16'b0101110110010011;    //sigmoid(1.000000) ≈ 0.731049
			6'b000011: sigmoid_out <= 16'b0110100010100110;    //sigmoid(1.500000) ≈ 0.817566
			6'b000100: sigmoid_out <= 16'b0111000010111110;    //sigmoid(2.000000) ≈ 0.880798
			6'b000101: sigmoid_out <= 16'b0111011001001010;    //sigmoid(2.500000) ≈ 0.924133
			6'b000110: sigmoid_out <= 16'b0111100111101110;    //sigmoid(3.000000) ≈ 0.952576
			6'b000111: sigmoid_out <= 16'b0111110000111111;    //sigmoid(3.500000) ≈ 0.970673
			6'b001000: sigmoid_out <= 16'b0111110110110011;    //sigmoid(4.000000) ≈ 0.982025
			6'b001001: sigmoid_out <= 16'b0111111010011000;    //sigmoid(4.500000) ≈ 0.989014
			6'b001010: sigmoid_out <= 16'b0111111100100101;    //sigmoid(5.000000) ≈ 0.993317
			6'b001011: sigmoid_out <= 16'b0111111101111011;    //sigmoid(5.500000) ≈ 0.995941
			6'b001100: sigmoid_out <= 16'b0111111110101111;    //sigmoid(6.000000) ≈ 0.997528
			6'b001101: sigmoid_out <= 16'b0111111111001111;    //sigmoid(6.500000) ≈ 0.998505
			6'b001110: sigmoid_out <= 16'b0111111111100010;    //sigmoid(7.000000) ≈ 0.999084
			6'b001111: sigmoid_out <= 16'b0111111111101110;    //sigmoid(7.500000) ≈ 0.999451
			6'b010000: sigmoid_out <= 16'b0111111111110101;    //sigmoid(8.000000) ≈ 0.999664
			6'b010001: sigmoid_out <= 16'b0111111111111001;    //sigmoid(8.500000) ≈ 0.999786
			6'b010010: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.000000) ≈ 0.999878
			6'b010011: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.500000) ≈ 0.999939
			6'b010100: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.000000) ≈ 0.999969
			6'b010101: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.500000) ≈ 0.999969
			6'b010110: sigmoid_out <= 16'b0111111111111111;    //sigmoid(11.000000) ≈ 0.999969
			6'b010111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.500000) ≈ 1.000000
			6'b011000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.000000) ≈ 1.000000
			6'b011001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.500000) ≈ 1.000000
			6'b011010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.000000) ≈ 1.000000
			6'b011011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.500000) ≈ 1.000000
			6'b011100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.000000) ≈ 1.000000
			6'b011101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.500000) ≈ 1.000000
			6'b011110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.000000) ≈ 1.000000
			6'b011111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.500000) ≈ 1.000000
			6'b100000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(16.000000) ≈ 1.000000
			6'b100001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(16.500000) ≈ 1.000000
			6'b100010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(17.000000) ≈ 1.000000
			6'b100011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(17.500000) ≈ 1.000000
			6'b100100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(18.000000) ≈ 1.000000
			6'b100101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(18.500000) ≈ 1.000000
			6'b100110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(19.000000) ≈ 1.000000
			6'b100111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(19.500000) ≈ 1.000000
			6'b101000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(20.000000) ≈ 1.000000
			6'b101001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(20.500000) ≈ 1.000000
			6'b101010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(21.000000) ≈ 1.000000
			6'b101011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(21.500000) ≈ 1.000000
			6'b101100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(22.000000) ≈ 1.000000
			6'b101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(22.500000) ≈ 1.000000
			6'b101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(23.000000) ≈ 1.000000
			6'b101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(23.500000) ≈ 1.000000
			6'b110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(24.000000) ≈ 1.000000
			6'b110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(24.500000) ≈ 1.000000
			6'b110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(25.000000) ≈ 1.000000
			6'b110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(25.500000) ≈ 1.000000
			6'b110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(26.000000) ≈ 1.000000
			6'b110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(26.500000) ≈ 1.000000
			6'b110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(27.000000) ≈ 1.000000
			6'b110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(27.500000) ≈ 1.000000
			6'b111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(28.000000) ≈ 1.000000
			6'b111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(28.500000) ≈ 1.000000
			6'b111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(29.000000) ≈ 1.000000
			6'b111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(29.500000) ≈ 1.000000
			6'b111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(30.000000) ≈ 1.000000
			6'b111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(30.500000) ≈ 1.000000
			6'b111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(31.000000) ≈ 1.000000
			6'b111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(31.500000) ≈ 1.000000

        endcase
    end
endmodule