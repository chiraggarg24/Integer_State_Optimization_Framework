//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2022-04-14 10:22:06.564762
// Design Name: vanilla
// Module Name: sigmoidLUT_in8b2p_out16b15p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 8 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in8b2p_out16b15p #(
    parameter PRECISION_INPUT_BITS = 8,
    parameter PRECISION_OUTPUT_BITS = 16
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			8'b00000000: sigmoid_out <= 16'b0100000000000000;    //sigmoid(0.000000) ≈ 0.500000
			8'b00000001: sigmoid_out <= 16'b0100011111110101;    //sigmoid(0.250000) ≈ 0.562164
			8'b00000010: sigmoid_out <= 16'b0100111110101101;    //sigmoid(0.500000) ≈ 0.622467
			8'b00000011: sigmoid_out <= 16'b0101011011101111;    //sigmoid(0.750000) ≈ 0.679169
			8'b00000100: sigmoid_out <= 16'b0101110110010011;    //sigmoid(1.000000) ≈ 0.731049
			8'b00000101: sigmoid_out <= 16'b0110001101111111;    //sigmoid(1.250000) ≈ 0.777313
			8'b00000110: sigmoid_out <= 16'b0110100010100110;    //sigmoid(1.500000) ≈ 0.817566
			8'b00000111: sigmoid_out <= 16'b0110110100001101;    //sigmoid(1.750000) ≈ 0.851959
			8'b00001000: sigmoid_out <= 16'b0111000010111110;    //sigmoid(2.000000) ≈ 0.880798
			8'b00001001: sigmoid_out <= 16'b0111001111001100;    //sigmoid(2.250000) ≈ 0.904663
			8'b00001010: sigmoid_out <= 16'b0111011001001010;    //sigmoid(2.500000) ≈ 0.924133
			8'b00001011: sigmoid_out <= 16'b0111100001001111;    //sigmoid(2.750000) ≈ 0.939911
			8'b00001100: sigmoid_out <= 16'b0111100111101110;    //sigmoid(3.000000) ≈ 0.952576
			8'b00001101: sigmoid_out <= 16'b0111101100111001;    //sigmoid(3.250000) ≈ 0.962677
			8'b00001110: sigmoid_out <= 16'b0111110000111111;    //sigmoid(3.500000) ≈ 0.970673
			8'b00001111: sigmoid_out <= 16'b0111110100001111;    //sigmoid(3.750000) ≈ 0.977020
			8'b00010000: sigmoid_out <= 16'b0111110110110011;    //sigmoid(4.000000) ≈ 0.982025
			8'b00010001: sigmoid_out <= 16'b0111111000110011;    //sigmoid(4.250000) ≈ 0.985931
			8'b00010010: sigmoid_out <= 16'b0111111010011000;    //sigmoid(4.500000) ≈ 0.989014
			8'b00010011: sigmoid_out <= 16'b0111111011100111;    //sigmoid(4.750000) ≈ 0.991425
			8'b00010100: sigmoid_out <= 16'b0111111100100101;    //sigmoid(5.000000) ≈ 0.993317
			8'b00010101: sigmoid_out <= 16'b0111111101010101;    //sigmoid(5.250000) ≈ 0.994781
			8'b00010110: sigmoid_out <= 16'b0111111101111011;    //sigmoid(5.500000) ≈ 0.995941
			8'b00010111: sigmoid_out <= 16'b0111111110011000;    //sigmoid(5.750000) ≈ 0.996826
			8'b00011000: sigmoid_out <= 16'b0111111110101111;    //sigmoid(6.000000) ≈ 0.997528
			8'b00011001: sigmoid_out <= 16'b0111111111000001;    //sigmoid(6.250000) ≈ 0.998077
			8'b00011010: sigmoid_out <= 16'b0111111111001111;    //sigmoid(6.500000) ≈ 0.998505
			8'b00011011: sigmoid_out <= 16'b0111111111011010;    //sigmoid(6.750000) ≈ 0.998840
			8'b00011100: sigmoid_out <= 16'b0111111111100010;    //sigmoid(7.000000) ≈ 0.999084
			8'b00011101: sigmoid_out <= 16'b0111111111101001;    //sigmoid(7.250000) ≈ 0.999298
			8'b00011110: sigmoid_out <= 16'b0111111111101110;    //sigmoid(7.500000) ≈ 0.999451
			8'b00011111: sigmoid_out <= 16'b0111111111110010;    //sigmoid(7.750000) ≈ 0.999573
			8'b00100000: sigmoid_out <= 16'b0111111111110101;    //sigmoid(8.000000) ≈ 0.999664
			8'b00100001: sigmoid_out <= 16'b0111111111110111;    //sigmoid(8.250000) ≈ 0.999725
			8'b00100010: sigmoid_out <= 16'b0111111111111001;    //sigmoid(8.500000) ≈ 0.999786
			8'b00100011: sigmoid_out <= 16'b0111111111111011;    //sigmoid(8.750000) ≈ 0.999847
			8'b00100100: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.000000) ≈ 0.999878
			8'b00100101: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.250000) ≈ 0.999908
			8'b00100110: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.500000) ≈ 0.999939
			8'b00100111: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.750000) ≈ 0.999939
			8'b00101000: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.000000) ≈ 0.999969
			8'b00101001: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.250000) ≈ 0.999969
			8'b00101010: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.500000) ≈ 0.999969
			8'b00101011: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.750000) ≈ 0.999969
			8'b00101100: sigmoid_out <= 16'b0111111111111111;    //sigmoid(11.000000) ≈ 0.999969
			8'b00101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.250000) ≈ 1.000000
			8'b00101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.500000) ≈ 1.000000
			8'b00101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.750000) ≈ 1.000000
			8'b00110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.000000) ≈ 1.000000
			8'b00110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.250000) ≈ 1.000000
			8'b00110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.500000) ≈ 1.000000
			8'b00110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.750000) ≈ 1.000000
			8'b00110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.000000) ≈ 1.000000
			8'b00110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.250000) ≈ 1.000000
			8'b00110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.500000) ≈ 1.000000
			8'b00110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.750000) ≈ 1.000000
			8'b00111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.000000) ≈ 1.000000
			8'b00111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.250000) ≈ 1.000000
			8'b00111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.500000) ≈ 1.000000
			8'b00111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.750000) ≈ 1.000000
			8'b00111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.000000) ≈ 1.000000
			8'b00111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.250000) ≈ 1.000000
			8'b00111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.500000) ≈ 1.000000
			8'b00111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.750000) ≈ 1.000000
			8'b01000000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(16.000000) ≈ 1.000000
			8'b01000001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(16.250000) ≈ 1.000000
			8'b01000010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(16.500000) ≈ 1.000000
			8'b01000011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(16.750000) ≈ 1.000000
			8'b01000100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(17.000000) ≈ 1.000000
			8'b01000101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(17.250000) ≈ 1.000000
			8'b01000110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(17.500000) ≈ 1.000000
			8'b01000111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(17.750000) ≈ 1.000000
			8'b01001000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(18.000000) ≈ 1.000000
			8'b01001001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(18.250000) ≈ 1.000000
			8'b01001010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(18.500000) ≈ 1.000000
			8'b01001011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(18.750000) ≈ 1.000000
			8'b01001100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(19.000000) ≈ 1.000000
			8'b01001101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(19.250000) ≈ 1.000000
			8'b01001110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(19.500000) ≈ 1.000000
			8'b01001111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(19.750000) ≈ 1.000000
			8'b01010000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(20.000000) ≈ 1.000000
			8'b01010001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(20.250000) ≈ 1.000000
			8'b01010010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(20.500000) ≈ 1.000000
			8'b01010011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(20.750000) ≈ 1.000000
			8'b01010100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(21.000000) ≈ 1.000000
			8'b01010101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(21.250000) ≈ 1.000000
			8'b01010110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(21.500000) ≈ 1.000000
			8'b01010111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(21.750000) ≈ 1.000000
			8'b01011000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(22.000000) ≈ 1.000000
			8'b01011001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(22.250000) ≈ 1.000000
			8'b01011010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(22.500000) ≈ 1.000000
			8'b01011011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(22.750000) ≈ 1.000000
			8'b01011100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(23.000000) ≈ 1.000000
			8'b01011101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(23.250000) ≈ 1.000000
			8'b01011110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(23.500000) ≈ 1.000000
			8'b01011111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(23.750000) ≈ 1.000000
			8'b01100000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(24.000000) ≈ 1.000000
			8'b01100001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(24.250000) ≈ 1.000000
			8'b01100010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(24.500000) ≈ 1.000000
			8'b01100011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(24.750000) ≈ 1.000000
			8'b01100100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(25.000000) ≈ 1.000000
			8'b01100101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(25.250000) ≈ 1.000000
			8'b01100110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(25.500000) ≈ 1.000000
			8'b01100111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(25.750000) ≈ 1.000000
			8'b01101000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(26.000000) ≈ 1.000000
			8'b01101001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(26.250000) ≈ 1.000000
			8'b01101010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(26.500000) ≈ 1.000000
			8'b01101011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(26.750000) ≈ 1.000000
			8'b01101100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(27.000000) ≈ 1.000000
			8'b01101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(27.250000) ≈ 1.000000
			8'b01101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(27.500000) ≈ 1.000000
			8'b01101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(27.750000) ≈ 1.000000
			8'b01110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(28.000000) ≈ 1.000000
			8'b01110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(28.250000) ≈ 1.000000
			8'b01110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(28.500000) ≈ 1.000000
			8'b01110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(28.750000) ≈ 1.000000
			8'b01110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(29.000000) ≈ 1.000000
			8'b01110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(29.250000) ≈ 1.000000
			8'b01110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(29.500000) ≈ 1.000000
			8'b01110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(29.750000) ≈ 1.000000
			8'b01111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(30.000000) ≈ 1.000000
			8'b01111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(30.250000) ≈ 1.000000
			8'b01111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(30.500000) ≈ 1.000000
			8'b01111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(30.750000) ≈ 1.000000
			8'b01111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(31.000000) ≈ 1.000000
			8'b01111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(31.250000) ≈ 1.000000
			8'b01111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(31.500000) ≈ 1.000000
			8'b01111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(31.750000) ≈ 1.000000
			8'b10000000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(32.000000) ≈ 1.000000
			8'b10000001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(32.250000) ≈ 1.000000
			8'b10000010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(32.500000) ≈ 1.000000
			8'b10000011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(32.750000) ≈ 1.000000
			8'b10000100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(33.000000) ≈ 1.000000
			8'b10000101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(33.250000) ≈ 1.000000
			8'b10000110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(33.500000) ≈ 1.000000
			8'b10000111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(33.750000) ≈ 1.000000
			8'b10001000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(34.000000) ≈ 1.000000
			8'b10001001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(34.250000) ≈ 1.000000
			8'b10001010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(34.500000) ≈ 1.000000
			8'b10001011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(34.750000) ≈ 1.000000
			8'b10001100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(35.000000) ≈ 1.000000
			8'b10001101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(35.250000) ≈ 1.000000
			8'b10001110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(35.500000) ≈ 1.000000
			8'b10001111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(35.750000) ≈ 1.000000
			8'b10010000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(36.000000) ≈ 1.000000
			8'b10010001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(36.250000) ≈ 1.000000
			8'b10010010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(36.500000) ≈ 1.000000
			8'b10010011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(36.750000) ≈ 1.000000
			8'b10010100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(37.000000) ≈ 1.000000
			8'b10010101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(37.250000) ≈ 1.000000
			8'b10010110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(37.500000) ≈ 1.000000
			8'b10010111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(37.750000) ≈ 1.000000
			8'b10011000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(38.000000) ≈ 1.000000
			8'b10011001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(38.250000) ≈ 1.000000
			8'b10011010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(38.500000) ≈ 1.000000
			8'b10011011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(38.750000) ≈ 1.000000
			8'b10011100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(39.000000) ≈ 1.000000
			8'b10011101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(39.250000) ≈ 1.000000
			8'b10011110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(39.500000) ≈ 1.000000
			8'b10011111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(39.750000) ≈ 1.000000
			8'b10100000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(40.000000) ≈ 1.000000
			8'b10100001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(40.250000) ≈ 1.000000
			8'b10100010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(40.500000) ≈ 1.000000
			8'b10100011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(40.750000) ≈ 1.000000
			8'b10100100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(41.000000) ≈ 1.000000
			8'b10100101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(41.250000) ≈ 1.000000
			8'b10100110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(41.500000) ≈ 1.000000
			8'b10100111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(41.750000) ≈ 1.000000
			8'b10101000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(42.000000) ≈ 1.000000
			8'b10101001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(42.250000) ≈ 1.000000
			8'b10101010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(42.500000) ≈ 1.000000
			8'b10101011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(42.750000) ≈ 1.000000
			8'b10101100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(43.000000) ≈ 1.000000
			8'b10101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(43.250000) ≈ 1.000000
			8'b10101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(43.500000) ≈ 1.000000
			8'b10101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(43.750000) ≈ 1.000000
			8'b10110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(44.000000) ≈ 1.000000
			8'b10110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(44.250000) ≈ 1.000000
			8'b10110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(44.500000) ≈ 1.000000
			8'b10110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(44.750000) ≈ 1.000000
			8'b10110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(45.000000) ≈ 1.000000
			8'b10110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(45.250000) ≈ 1.000000
			8'b10110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(45.500000) ≈ 1.000000
			8'b10110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(45.750000) ≈ 1.000000
			8'b10111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(46.000000) ≈ 1.000000
			8'b10111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(46.250000) ≈ 1.000000
			8'b10111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(46.500000) ≈ 1.000000
			8'b10111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(46.750000) ≈ 1.000000
			8'b10111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(47.000000) ≈ 1.000000
			8'b10111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(47.250000) ≈ 1.000000
			8'b10111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(47.500000) ≈ 1.000000
			8'b10111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(47.750000) ≈ 1.000000
			8'b11000000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(48.000000) ≈ 1.000000
			8'b11000001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(48.250000) ≈ 1.000000
			8'b11000010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(48.500000) ≈ 1.000000
			8'b11000011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(48.750000) ≈ 1.000000
			8'b11000100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(49.000000) ≈ 1.000000
			8'b11000101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(49.250000) ≈ 1.000000
			8'b11000110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(49.500000) ≈ 1.000000
			8'b11000111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(49.750000) ≈ 1.000000
			8'b11001000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(50.000000) ≈ 1.000000
			8'b11001001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(50.250000) ≈ 1.000000
			8'b11001010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(50.500000) ≈ 1.000000
			8'b11001011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(50.750000) ≈ 1.000000
			8'b11001100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(51.000000) ≈ 1.000000
			8'b11001101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(51.250000) ≈ 1.000000
			8'b11001110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(51.500000) ≈ 1.000000
			8'b11001111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(51.750000) ≈ 1.000000
			8'b11010000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(52.000000) ≈ 1.000000
			8'b11010001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(52.250000) ≈ 1.000000
			8'b11010010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(52.500000) ≈ 1.000000
			8'b11010011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(52.750000) ≈ 1.000000
			8'b11010100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(53.000000) ≈ 1.000000
			8'b11010101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(53.250000) ≈ 1.000000
			8'b11010110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(53.500000) ≈ 1.000000
			8'b11010111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(53.750000) ≈ 1.000000
			8'b11011000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(54.000000) ≈ 1.000000
			8'b11011001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(54.250000) ≈ 1.000000
			8'b11011010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(54.500000) ≈ 1.000000
			8'b11011011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(54.750000) ≈ 1.000000
			8'b11011100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(55.000000) ≈ 1.000000
			8'b11011101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(55.250000) ≈ 1.000000
			8'b11011110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(55.500000) ≈ 1.000000
			8'b11011111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(55.750000) ≈ 1.000000
			8'b11100000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(56.000000) ≈ 1.000000
			8'b11100001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(56.250000) ≈ 1.000000
			8'b11100010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(56.500000) ≈ 1.000000
			8'b11100011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(56.750000) ≈ 1.000000
			8'b11100100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(57.000000) ≈ 1.000000
			8'b11100101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(57.250000) ≈ 1.000000
			8'b11100110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(57.500000) ≈ 1.000000
			8'b11100111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(57.750000) ≈ 1.000000
			8'b11101000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(58.000000) ≈ 1.000000
			8'b11101001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(58.250000) ≈ 1.000000
			8'b11101010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(58.500000) ≈ 1.000000
			8'b11101011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(58.750000) ≈ 1.000000
			8'b11101100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(59.000000) ≈ 1.000000
			8'b11101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(59.250000) ≈ 1.000000
			8'b11101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(59.500000) ≈ 1.000000
			8'b11101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(59.750000) ≈ 1.000000
			8'b11110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(60.000000) ≈ 1.000000
			8'b11110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(60.250000) ≈ 1.000000
			8'b11110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(60.500000) ≈ 1.000000
			8'b11110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(60.750000) ≈ 1.000000
			8'b11110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(61.000000) ≈ 1.000000
			8'b11110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(61.250000) ≈ 1.000000
			8'b11110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(61.500000) ≈ 1.000000
			8'b11110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(61.750000) ≈ 1.000000
			8'b11111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(62.000000) ≈ 1.000000
			8'b11111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(62.250000) ≈ 1.000000
			8'b11111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(62.500000) ≈ 1.000000
			8'b11111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(62.750000) ≈ 1.000000
			8'b11111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(63.000000) ≈ 1.000000
			8'b11111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(63.250000) ≈ 1.000000
			8'b11111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(63.500000) ≈ 1.000000
			8'b11111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(63.750000) ≈ 1.000000

        endcase
    end
endmodule