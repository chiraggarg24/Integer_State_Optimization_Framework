//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2022-06-23 15:11:55.058043
// Design Name: vanilla
// Module Name: sigmoidLUT_in7b3p_out16b15p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 7 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in7b3p_out16b15p #(
    parameter PRECISION_INPUT_BITS = 7,
    parameter PRECISION_OUTPUT_BITS = 16
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			7'b0000000: sigmoid_out <= 16'b0100000000000000;    //sigmoid(0.000000) ≈ 0.500000
			7'b0000001: sigmoid_out <= 16'b0100001111111111;    //sigmoid(0.125000) ≈ 0.531219
			7'b0000010: sigmoid_out <= 16'b0100011111110101;    //sigmoid(0.250000) ≈ 0.562164
			7'b0000011: sigmoid_out <= 16'b0100101111011100;    //sigmoid(0.375000) ≈ 0.592651
			7'b0000100: sigmoid_out <= 16'b0100111110101101;    //sigmoid(0.500000) ≈ 0.622467
			7'b0000101: sigmoid_out <= 16'b0101001101100000;    //sigmoid(0.625000) ≈ 0.651367
			7'b0000110: sigmoid_out <= 16'b0101011011101111;    //sigmoid(0.750000) ≈ 0.679169
			7'b0000111: sigmoid_out <= 16'b0101101001010111;    //sigmoid(0.875000) ≈ 0.705780
			7'b0001000: sigmoid_out <= 16'b0101110110010011;    //sigmoid(1.000000) ≈ 0.731049
			7'b0001001: sigmoid_out <= 16'b0110000010100001;    //sigmoid(1.125000) ≈ 0.754913
			7'b0001010: sigmoid_out <= 16'b0110001101111111;    //sigmoid(1.250000) ≈ 0.777313
			7'b0001011: sigmoid_out <= 16'b0110011000101011;    //sigmoid(1.375000) ≈ 0.798187
			7'b0001100: sigmoid_out <= 16'b0110100010100110;    //sigmoid(1.500000) ≈ 0.817566
			7'b0001101: sigmoid_out <= 16'b0110101011110001;    //sigmoid(1.625000) ≈ 0.835480
			7'b0001110: sigmoid_out <= 16'b0110110100001101;    //sigmoid(1.750000) ≈ 0.851959
			7'b0001111: sigmoid_out <= 16'b0110111011111011;    //sigmoid(1.875000) ≈ 0.867035
			7'b0010000: sigmoid_out <= 16'b0111000010111110;    //sigmoid(2.000000) ≈ 0.880798
			7'b0010001: sigmoid_out <= 16'b0111001001011000;    //sigmoid(2.125000) ≈ 0.893311
			7'b0010010: sigmoid_out <= 16'b0111001111001100;    //sigmoid(2.250000) ≈ 0.904663
			7'b0010011: sigmoid_out <= 16'b0111010100011011;    //sigmoid(2.375000) ≈ 0.914886
			7'b0010100: sigmoid_out <= 16'b0111011001001010;    //sigmoid(2.500000) ≈ 0.924133
			7'b0010101: sigmoid_out <= 16'b0111011101011011;    //sigmoid(2.625000) ≈ 0.932465
			7'b0010110: sigmoid_out <= 16'b0111100001001111;    //sigmoid(2.750000) ≈ 0.939911
			7'b0010111: sigmoid_out <= 16'b0111100100101010;    //sigmoid(2.875000) ≈ 0.946594
			7'b0011000: sigmoid_out <= 16'b0111100111101110;    //sigmoid(3.000000) ≈ 0.952576
			7'b0011001: sigmoid_out <= 16'b0111101010011101;    //sigmoid(3.125000) ≈ 0.957916
			7'b0011010: sigmoid_out <= 16'b0111101100111001;    //sigmoid(3.250000) ≈ 0.962677
			7'b0011011: sigmoid_out <= 16'b0111101111000100;    //sigmoid(3.375000) ≈ 0.966919
			7'b0011100: sigmoid_out <= 16'b0111110000111111;    //sigmoid(3.500000) ≈ 0.970673
			7'b0011101: sigmoid_out <= 16'b0111110010101101;    //sigmoid(3.625000) ≈ 0.974030
			7'b0011110: sigmoid_out <= 16'b0111110100001111;    //sigmoid(3.750000) ≈ 0.977020
			7'b0011111: sigmoid_out <= 16'b0111110101100110;    //sigmoid(3.875000) ≈ 0.979675
			7'b0100000: sigmoid_out <= 16'b0111110110110011;    //sigmoid(4.000000) ≈ 0.982025
			7'b0100001: sigmoid_out <= 16'b0111110111110111;    //sigmoid(4.125000) ≈ 0.984100
			7'b0100010: sigmoid_out <= 16'b0111111000110011;    //sigmoid(4.250000) ≈ 0.985931
			7'b0100011: sigmoid_out <= 16'b0111111001101001;    //sigmoid(4.375000) ≈ 0.987579
			7'b0100100: sigmoid_out <= 16'b0111111010011000;    //sigmoid(4.500000) ≈ 0.989014
			7'b0100101: sigmoid_out <= 16'b0111111011000010;    //sigmoid(4.625000) ≈ 0.990295
			7'b0100110: sigmoid_out <= 16'b0111111011100111;    //sigmoid(4.750000) ≈ 0.991425
			7'b0100111: sigmoid_out <= 16'b0111111100001000;    //sigmoid(4.875000) ≈ 0.992432
			7'b0101000: sigmoid_out <= 16'b0111111100100101;    //sigmoid(5.000000) ≈ 0.993317
			7'b0101001: sigmoid_out <= 16'b0111111100111110;    //sigmoid(5.125000) ≈ 0.994080
			7'b0101010: sigmoid_out <= 16'b0111111101010101;    //sigmoid(5.250000) ≈ 0.994781
			7'b0101011: sigmoid_out <= 16'b0111111101101001;    //sigmoid(5.375000) ≈ 0.995392
			7'b0101100: sigmoid_out <= 16'b0111111101111011;    //sigmoid(5.500000) ≈ 0.995941
			7'b0101101: sigmoid_out <= 16'b0111111110001010;    //sigmoid(5.625000) ≈ 0.996399
			7'b0101110: sigmoid_out <= 16'b0111111110011000;    //sigmoid(5.750000) ≈ 0.996826
			7'b0101111: sigmoid_out <= 16'b0111111110100100;    //sigmoid(5.875000) ≈ 0.997192
			7'b0110000: sigmoid_out <= 16'b0111111110101111;    //sigmoid(6.000000) ≈ 0.997528
			7'b0110001: sigmoid_out <= 16'b0111111110111000;    //sigmoid(6.125000) ≈ 0.997803
			7'b0110010: sigmoid_out <= 16'b0111111111000001;    //sigmoid(6.250000) ≈ 0.998077
			7'b0110011: sigmoid_out <= 16'b0111111111001000;    //sigmoid(6.375000) ≈ 0.998291
			7'b0110100: sigmoid_out <= 16'b0111111111001111;    //sigmoid(6.500000) ≈ 0.998505
			7'b0110101: sigmoid_out <= 16'b0111111111010101;    //sigmoid(6.625000) ≈ 0.998688
			7'b0110110: sigmoid_out <= 16'b0111111111011010;    //sigmoid(6.750000) ≈ 0.998840
			7'b0110111: sigmoid_out <= 16'b0111111111011110;    //sigmoid(6.875000) ≈ 0.998962
			7'b0111000: sigmoid_out <= 16'b0111111111100010;    //sigmoid(7.000000) ≈ 0.999084
			7'b0111001: sigmoid_out <= 16'b0111111111100110;    //sigmoid(7.125000) ≈ 0.999207
			7'b0111010: sigmoid_out <= 16'b0111111111101001;    //sigmoid(7.250000) ≈ 0.999298
			7'b0111011: sigmoid_out <= 16'b0111111111101011;    //sigmoid(7.375000) ≈ 0.999359
			7'b0111100: sigmoid_out <= 16'b0111111111101110;    //sigmoid(7.500000) ≈ 0.999451
			7'b0111101: sigmoid_out <= 16'b0111111111110000;    //sigmoid(7.625000) ≈ 0.999512
			7'b0111110: sigmoid_out <= 16'b0111111111110010;    //sigmoid(7.750000) ≈ 0.999573
			7'b0111111: sigmoid_out <= 16'b0111111111110100;    //sigmoid(7.875000) ≈ 0.999634
			7'b1000000: sigmoid_out <= 16'b0111111111110101;    //sigmoid(8.000000) ≈ 0.999664
			7'b1000001: sigmoid_out <= 16'b0111111111110110;    //sigmoid(8.125000) ≈ 0.999695
			7'b1000010: sigmoid_out <= 16'b0111111111110111;    //sigmoid(8.250000) ≈ 0.999725
			7'b1000011: sigmoid_out <= 16'b0111111111111000;    //sigmoid(8.375000) ≈ 0.999756
			7'b1000100: sigmoid_out <= 16'b0111111111111001;    //sigmoid(8.500000) ≈ 0.999786
			7'b1000101: sigmoid_out <= 16'b0111111111111010;    //sigmoid(8.625000) ≈ 0.999817
			7'b1000110: sigmoid_out <= 16'b0111111111111011;    //sigmoid(8.750000) ≈ 0.999847
			7'b1000111: sigmoid_out <= 16'b0111111111111011;    //sigmoid(8.875000) ≈ 0.999847
			7'b1001000: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.000000) ≈ 0.999878
			7'b1001001: sigmoid_out <= 16'b0111111111111100;    //sigmoid(9.125000) ≈ 0.999878
			7'b1001010: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.250000) ≈ 0.999908
			7'b1001011: sigmoid_out <= 16'b0111111111111101;    //sigmoid(9.375000) ≈ 0.999908
			7'b1001100: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.500000) ≈ 0.999939
			7'b1001101: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.625000) ≈ 0.999939
			7'b1001110: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.750000) ≈ 0.999939
			7'b1001111: sigmoid_out <= 16'b0111111111111110;    //sigmoid(9.875000) ≈ 0.999939
			7'b1010000: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.000000) ≈ 0.999969
			7'b1010001: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.125000) ≈ 0.999969
			7'b1010010: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.250000) ≈ 0.999969
			7'b1010011: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.375000) ≈ 0.999969
			7'b1010100: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.500000) ≈ 0.999969
			7'b1010101: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.625000) ≈ 0.999969
			7'b1010110: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.750000) ≈ 0.999969
			7'b1010111: sigmoid_out <= 16'b0111111111111111;    //sigmoid(10.875000) ≈ 0.999969
			7'b1011000: sigmoid_out <= 16'b0111111111111111;    //sigmoid(11.000000) ≈ 0.999969
			7'b1011001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.125000) ≈ 1.000000
			7'b1011010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.250000) ≈ 1.000000
			7'b1011011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.375000) ≈ 1.000000
			7'b1011100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.500000) ≈ 1.000000
			7'b1011101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.625000) ≈ 1.000000
			7'b1011110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.750000) ≈ 1.000000
			7'b1011111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(11.875000) ≈ 1.000000
			7'b1100000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.000000) ≈ 1.000000
			7'b1100001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.125000) ≈ 1.000000
			7'b1100010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.250000) ≈ 1.000000
			7'b1100011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.375000) ≈ 1.000000
			7'b1100100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.500000) ≈ 1.000000
			7'b1100101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.625000) ≈ 1.000000
			7'b1100110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.750000) ≈ 1.000000
			7'b1100111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(12.875000) ≈ 1.000000
			7'b1101000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.000000) ≈ 1.000000
			7'b1101001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.125000) ≈ 1.000000
			7'b1101010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.250000) ≈ 1.000000
			7'b1101011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.375000) ≈ 1.000000
			7'b1101100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.500000) ≈ 1.000000
			7'b1101101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.625000) ≈ 1.000000
			7'b1101110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.750000) ≈ 1.000000
			7'b1101111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(13.875000) ≈ 1.000000
			7'b1110000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.000000) ≈ 1.000000
			7'b1110001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.125000) ≈ 1.000000
			7'b1110010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.250000) ≈ 1.000000
			7'b1110011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.375000) ≈ 1.000000
			7'b1110100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.500000) ≈ 1.000000
			7'b1110101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.625000) ≈ 1.000000
			7'b1110110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.750000) ≈ 1.000000
			7'b1110111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(14.875000) ≈ 1.000000
			7'b1111000: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.000000) ≈ 1.000000
			7'b1111001: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.125000) ≈ 1.000000
			7'b1111010: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.250000) ≈ 1.000000
			7'b1111011: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.375000) ≈ 1.000000
			7'b1111100: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.500000) ≈ 1.000000
			7'b1111101: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.625000) ≈ 1.000000
			7'b1111110: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.750000) ≈ 1.000000
			7'b1111111: sigmoid_out <= 16'b1000000000000000;    //sigmoid(15.875000) ≈ 1.000000

        endcase
    end
endmodule