//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-06-28 15:12:04.368345
// Design Name: vanilla
// Module Name: sigmoidLUT_in7b4p_out10b10p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 7 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in7b4p_out10b10p #(
    parameter PRECISION_INPUT_BITS = 7,
    parameter PRECISION_OUTPUT_BITS = 10
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			7'b0000000: sigmoid_out <= 10'b1000000000;    //sigmoid(0.000000) ≈ 0.500000
			7'b0000001: sigmoid_out <= 10'b1000010000;    //sigmoid(0.062500) ≈ 0.515625
			7'b0000010: sigmoid_out <= 10'b1000100000;    //sigmoid(0.125000) ≈ 0.531250
			7'b0000011: sigmoid_out <= 10'b1000110000;    //sigmoid(0.187500) ≈ 0.546875
			7'b0000100: sigmoid_out <= 10'b1001000000;    //sigmoid(0.250000) ≈ 0.562500
			7'b0000101: sigmoid_out <= 10'b1001001111;    //sigmoid(0.312500) ≈ 0.577148
			7'b0000110: sigmoid_out <= 10'b1001011111;    //sigmoid(0.375000) ≈ 0.592773
			7'b0000111: sigmoid_out <= 10'b1001101110;    //sigmoid(0.437500) ≈ 0.607422
			7'b0001000: sigmoid_out <= 10'b1001111101;    //sigmoid(0.500000) ≈ 0.622070
			7'b0001001: sigmoid_out <= 10'b1010001100;    //sigmoid(0.562500) ≈ 0.636719
			7'b0001010: sigmoid_out <= 10'b1010011011;    //sigmoid(0.625000) ≈ 0.651367
			7'b0001011: sigmoid_out <= 10'b1010101001;    //sigmoid(0.687500) ≈ 0.665039
			7'b0001100: sigmoid_out <= 10'b1010110111;    //sigmoid(0.750000) ≈ 0.678711
			7'b0001101: sigmoid_out <= 10'b1011000101;    //sigmoid(0.812500) ≈ 0.692383
			7'b0001110: sigmoid_out <= 10'b1011010011;    //sigmoid(0.875000) ≈ 0.706055
			7'b0001111: sigmoid_out <= 10'b1011100000;    //sigmoid(0.937500) ≈ 0.718750
			7'b0010000: sigmoid_out <= 10'b1011101101;    //sigmoid(1.000000) ≈ 0.731445
			7'b0010001: sigmoid_out <= 10'b1011111001;    //sigmoid(1.062500) ≈ 0.743164
			7'b0010010: sigmoid_out <= 10'b1100000101;    //sigmoid(1.125000) ≈ 0.754883
			7'b0010011: sigmoid_out <= 10'b1100010001;    //sigmoid(1.187500) ≈ 0.766602
			7'b0010100: sigmoid_out <= 10'b1100011100;    //sigmoid(1.250000) ≈ 0.777344
			7'b0010101: sigmoid_out <= 10'b1100100111;    //sigmoid(1.312500) ≈ 0.788086
			7'b0010110: sigmoid_out <= 10'b1100110001;    //sigmoid(1.375000) ≈ 0.797852
			7'b0010111: sigmoid_out <= 10'b1100111011;    //sigmoid(1.437500) ≈ 0.807617
			7'b0011000: sigmoid_out <= 10'b1101000101;    //sigmoid(1.500000) ≈ 0.817383
			7'b0011001: sigmoid_out <= 10'b1101001111;    //sigmoid(1.562500) ≈ 0.827148
			7'b0011010: sigmoid_out <= 10'b1101011000;    //sigmoid(1.625000) ≈ 0.835938
			7'b0011011: sigmoid_out <= 10'b1101100000;    //sigmoid(1.687500) ≈ 0.843750
			7'b0011100: sigmoid_out <= 10'b1101101000;    //sigmoid(1.750000) ≈ 0.851562
			7'b0011101: sigmoid_out <= 10'b1101110000;    //sigmoid(1.812500) ≈ 0.859375
			7'b0011110: sigmoid_out <= 10'b1101111000;    //sigmoid(1.875000) ≈ 0.867188
			7'b0011111: sigmoid_out <= 10'b1101111111;    //sigmoid(1.937500) ≈ 0.874023
			7'b0100000: sigmoid_out <= 10'b1110000110;    //sigmoid(2.000000) ≈ 0.880859
			7'b0100001: sigmoid_out <= 10'b1110001100;    //sigmoid(2.062500) ≈ 0.886719
			7'b0100010: sigmoid_out <= 10'b1110010011;    //sigmoid(2.125000) ≈ 0.893555
			7'b0100011: sigmoid_out <= 10'b1110011001;    //sigmoid(2.187500) ≈ 0.899414
			7'b0100100: sigmoid_out <= 10'b1110011110;    //sigmoid(2.250000) ≈ 0.904297
			7'b0100101: sigmoid_out <= 10'b1110100100;    //sigmoid(2.312500) ≈ 0.910156
			7'b0100110: sigmoid_out <= 10'b1110101001;    //sigmoid(2.375000) ≈ 0.915039
			7'b0100111: sigmoid_out <= 10'b1110101110;    //sigmoid(2.437500) ≈ 0.919922
			7'b0101000: sigmoid_out <= 10'b1110110010;    //sigmoid(2.500000) ≈ 0.923828
			7'b0101001: sigmoid_out <= 10'b1110110111;    //sigmoid(2.562500) ≈ 0.928711
			7'b0101010: sigmoid_out <= 10'b1110111011;    //sigmoid(2.625000) ≈ 0.932617
			7'b0101011: sigmoid_out <= 10'b1110111111;    //sigmoid(2.687500) ≈ 0.936523
			7'b0101100: sigmoid_out <= 10'b1111000010;    //sigmoid(2.750000) ≈ 0.939453
			7'b0101101: sigmoid_out <= 10'b1111000110;    //sigmoid(2.812500) ≈ 0.943359
			7'b0101110: sigmoid_out <= 10'b1111001001;    //sigmoid(2.875000) ≈ 0.946289
			7'b0101111: sigmoid_out <= 10'b1111001100;    //sigmoid(2.937500) ≈ 0.949219
			7'b0110000: sigmoid_out <= 10'b1111001111;    //sigmoid(3.000000) ≈ 0.952148
			7'b0110001: sigmoid_out <= 10'b1111010010;    //sigmoid(3.062500) ≈ 0.955078
			7'b0110010: sigmoid_out <= 10'b1111010101;    //sigmoid(3.125000) ≈ 0.958008
			7'b0110011: sigmoid_out <= 10'b1111010111;    //sigmoid(3.187500) ≈ 0.959961
			7'b0110100: sigmoid_out <= 10'b1111011010;    //sigmoid(3.250000) ≈ 0.962891
			7'b0110101: sigmoid_out <= 10'b1111011100;    //sigmoid(3.312500) ≈ 0.964844
			7'b0110110: sigmoid_out <= 10'b1111011110;    //sigmoid(3.375000) ≈ 0.966797
			7'b0110111: sigmoid_out <= 10'b1111100000;    //sigmoid(3.437500) ≈ 0.968750
			7'b0111000: sigmoid_out <= 10'b1111100010;    //sigmoid(3.500000) ≈ 0.970703
			7'b0111001: sigmoid_out <= 10'b1111100100;    //sigmoid(3.562500) ≈ 0.972656
			7'b0111010: sigmoid_out <= 10'b1111100101;    //sigmoid(3.625000) ≈ 0.973633
			7'b0111011: sigmoid_out <= 10'b1111100111;    //sigmoid(3.687500) ≈ 0.975586
			7'b0111100: sigmoid_out <= 10'b1111101000;    //sigmoid(3.750000) ≈ 0.976562
			7'b0111101: sigmoid_out <= 10'b1111101010;    //sigmoid(3.812500) ≈ 0.978516
			7'b0111110: sigmoid_out <= 10'b1111101011;    //sigmoid(3.875000) ≈ 0.979492
			7'b0111111: sigmoid_out <= 10'b1111101100;    //sigmoid(3.937500) ≈ 0.980469
			7'b1000000: sigmoid_out <= 10'b1111101110;    //sigmoid(4.000000) ≈ 0.982422
			7'b1000001: sigmoid_out <= 10'b1111101111;    //sigmoid(4.062500) ≈ 0.983398
			7'b1000010: sigmoid_out <= 10'b1111110000;    //sigmoid(4.125000) ≈ 0.984375
			7'b1000011: sigmoid_out <= 10'b1111110001;    //sigmoid(4.187500) ≈ 0.985352
			7'b1000100: sigmoid_out <= 10'b1111110010;    //sigmoid(4.250000) ≈ 0.986328
			7'b1000101: sigmoid_out <= 10'b1111110010;    //sigmoid(4.312500) ≈ 0.986328
			7'b1000110: sigmoid_out <= 10'b1111110011;    //sigmoid(4.375000) ≈ 0.987305
			7'b1000111: sigmoid_out <= 10'b1111110100;    //sigmoid(4.437500) ≈ 0.988281
			7'b1001000: sigmoid_out <= 10'b1111110101;    //sigmoid(4.500000) ≈ 0.989258
			7'b1001001: sigmoid_out <= 10'b1111110101;    //sigmoid(4.562500) ≈ 0.989258
			7'b1001010: sigmoid_out <= 10'b1111110110;    //sigmoid(4.625000) ≈ 0.990234
			7'b1001011: sigmoid_out <= 10'b1111110111;    //sigmoid(4.687500) ≈ 0.991211
			7'b1001100: sigmoid_out <= 10'b1111110111;    //sigmoid(4.750000) ≈ 0.991211
			7'b1001101: sigmoid_out <= 10'b1111111000;    //sigmoid(4.812500) ≈ 0.992188
			7'b1001110: sigmoid_out <= 10'b1111111000;    //sigmoid(4.875000) ≈ 0.992188
			7'b1001111: sigmoid_out <= 10'b1111111001;    //sigmoid(4.937500) ≈ 0.993164
			7'b1010000: sigmoid_out <= 10'b1111111001;    //sigmoid(5.000000) ≈ 0.993164
			7'b1010001: sigmoid_out <= 10'b1111111010;    //sigmoid(5.062500) ≈ 0.994141
			7'b1010010: sigmoid_out <= 10'b1111111010;    //sigmoid(5.125000) ≈ 0.994141
			7'b1010011: sigmoid_out <= 10'b1111111010;    //sigmoid(5.187500) ≈ 0.994141
			7'b1010100: sigmoid_out <= 10'b1111111011;    //sigmoid(5.250000) ≈ 0.995117
			7'b1010101: sigmoid_out <= 10'b1111111011;    //sigmoid(5.312500) ≈ 0.995117
			7'b1010110: sigmoid_out <= 10'b1111111011;    //sigmoid(5.375000) ≈ 0.995117
			7'b1010111: sigmoid_out <= 10'b1111111100;    //sigmoid(5.437500) ≈ 0.996094
			7'b1011000: sigmoid_out <= 10'b1111111100;    //sigmoid(5.500000) ≈ 0.996094
			7'b1011001: sigmoid_out <= 10'b1111111100;    //sigmoid(5.562500) ≈ 0.996094
			7'b1011010: sigmoid_out <= 10'b1111111100;    //sigmoid(5.625000) ≈ 0.996094
			7'b1011011: sigmoid_out <= 10'b1111111101;    //sigmoid(5.687500) ≈ 0.997070
			7'b1011100: sigmoid_out <= 10'b1111111101;    //sigmoid(5.750000) ≈ 0.997070
			7'b1011101: sigmoid_out <= 10'b1111111101;    //sigmoid(5.812500) ≈ 0.997070
			7'b1011110: sigmoid_out <= 10'b1111111101;    //sigmoid(5.875000) ≈ 0.997070
			7'b1011111: sigmoid_out <= 10'b1111111101;    //sigmoid(5.937500) ≈ 0.997070
			7'b1100000: sigmoid_out <= 10'b1111111101;    //sigmoid(6.000000) ≈ 0.997070
			7'b1100001: sigmoid_out <= 10'b1111111110;    //sigmoid(6.062500) ≈ 0.998047
			7'b1100010: sigmoid_out <= 10'b1111111110;    //sigmoid(6.125000) ≈ 0.998047
			7'b1100011: sigmoid_out <= 10'b1111111110;    //sigmoid(6.187500) ≈ 0.998047
			7'b1100100: sigmoid_out <= 10'b1111111110;    //sigmoid(6.250000) ≈ 0.998047
			7'b1100101: sigmoid_out <= 10'b1111111110;    //sigmoid(6.312500) ≈ 0.998047
			7'b1100110: sigmoid_out <= 10'b1111111110;    //sigmoid(6.375000) ≈ 0.998047
			7'b1100111: sigmoid_out <= 10'b1111111110;    //sigmoid(6.437500) ≈ 0.998047
			7'b1101000: sigmoid_out <= 10'b1111111110;    //sigmoid(6.500000) ≈ 0.998047
			7'b1101001: sigmoid_out <= 10'b1111111111;    //sigmoid(6.562500) ≈ 0.999023
			7'b1101010: sigmoid_out <= 10'b1111111111;    //sigmoid(6.625000) ≈ 0.999023
			7'b1101011: sigmoid_out <= 10'b1111111111;    //sigmoid(6.687500) ≈ 0.999023
			7'b1101100: sigmoid_out <= 10'b1111111111;    //sigmoid(6.750000) ≈ 0.999023
			7'b1101101: sigmoid_out <= 10'b1111111111;    //sigmoid(6.812500) ≈ 0.999023
			7'b1101110: sigmoid_out <= 10'b1111111111;    //sigmoid(6.875000) ≈ 0.999023
			7'b1101111: sigmoid_out <= 10'b1111111111;    //sigmoid(6.937500) ≈ 0.999023
			7'b1110000: sigmoid_out <= 10'b1111111111;    //sigmoid(7.000000) ≈ 0.999023
			7'b1110001: sigmoid_out <= 10'b1111111111;    //sigmoid(7.062500) ≈ 0.999023
			7'b1110010: sigmoid_out <= 10'b1111111111;    //sigmoid(7.125000) ≈ 0.999023
			7'b1110011: sigmoid_out <= 10'b1111111111;    //sigmoid(7.187500) ≈ 0.999023
			7'b1110100: sigmoid_out <= 10'b1111111111;    //sigmoid(7.250000) ≈ 0.999023
			7'b1110101: sigmoid_out <= 10'b1111111111;    //sigmoid(7.312500) ≈ 0.999023
			7'b1110110: sigmoid_out <= 10'b1111111111;    //sigmoid(7.375000) ≈ 0.999023
			7'b1110111: sigmoid_out <= 10'b1111111111;    //sigmoid(7.437500) ≈ 0.999023
			7'b1111000: sigmoid_out <= 10'b1111111111;    //sigmoid(7.500000) ≈ 0.999023
			7'b1111001: sigmoid_out <= 10'b1111111111;    //sigmoid(7.562500) ≈ 0.999023
			7'b1111010: sigmoid_out <= 10'b1111111111;    //sigmoid(7.625000) ≈ 0.999023
			7'b1111011: sigmoid_out <= 10'b1111111111;    //sigmoid(7.687500) ≈ 0.999023
			7'b1111100: sigmoid_out <= 10'b1111111111;    //sigmoid(7.750000) ≈ 0.999023
			7'b1111101: sigmoid_out <= 10'b1111111111;    //sigmoid(7.812500) ≈ 0.999023
			7'b1111110: sigmoid_out <= 10'b1111111111;    //sigmoid(7.875000) ≈ 0.999023
			7'b1111111: sigmoid_out <= 10'b1111111111;    //sigmoid(7.937500) ≈ 0.999023

        endcase
    end
endmodule