//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
// 
// Create Date: 2019-06-28 11:49:47.978804
// Design Name: vanilla
// Module Name: sigmoidLUT_7bit_4point
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 7 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
// 
// Additional Comments: Generated by LUT_generator_sigmoid.py
// 
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_7bit_4point #(
    parameter PRECISION_BITS = 7
)(
    input[PRECISION_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			7'b0000000: sigmoid_out <= 7'b0001000;    //sigmoid(0.000000) ≈ 0.500000
			7'b0000001: sigmoid_out <= 7'b0001000;    //sigmoid(0.062500) ≈ 0.500000
			7'b0000010: sigmoid_out <= 7'b0001000;    //sigmoid(0.125000) ≈ 0.500000
			7'b0000011: sigmoid_out <= 7'b0001001;    //sigmoid(0.187500) ≈ 0.562500
			7'b0000100: sigmoid_out <= 7'b0001001;    //sigmoid(0.250000) ≈ 0.562500
			7'b0000101: sigmoid_out <= 7'b0001001;    //sigmoid(0.312500) ≈ 0.562500
			7'b0000110: sigmoid_out <= 7'b0001001;    //sigmoid(0.375000) ≈ 0.562500
			7'b0000111: sigmoid_out <= 7'b0001010;    //sigmoid(0.437500) ≈ 0.625000
			7'b0001000: sigmoid_out <= 7'b0001010;    //sigmoid(0.500000) ≈ 0.625000
			7'b0001001: sigmoid_out <= 7'b0001010;    //sigmoid(0.562500) ≈ 0.625000
			7'b0001010: sigmoid_out <= 7'b0001010;    //sigmoid(0.625000) ≈ 0.625000
			7'b0001011: sigmoid_out <= 7'b0001011;    //sigmoid(0.687500) ≈ 0.687500
			7'b0001100: sigmoid_out <= 7'b0001011;    //sigmoid(0.750000) ≈ 0.687500
			7'b0001101: sigmoid_out <= 7'b0001011;    //sigmoid(0.812500) ≈ 0.687500
			7'b0001110: sigmoid_out <= 7'b0001011;    //sigmoid(0.875000) ≈ 0.687500
			7'b0001111: sigmoid_out <= 7'b0001011;    //sigmoid(0.937500) ≈ 0.687500
			7'b0010000: sigmoid_out <= 7'b0001100;    //sigmoid(1.000000) ≈ 0.750000
			7'b0010001: sigmoid_out <= 7'b0001100;    //sigmoid(1.062500) ≈ 0.750000
			7'b0010010: sigmoid_out <= 7'b0001100;    //sigmoid(1.125000) ≈ 0.750000
			7'b0010011: sigmoid_out <= 7'b0001100;    //sigmoid(1.187500) ≈ 0.750000
			7'b0010100: sigmoid_out <= 7'b0001100;    //sigmoid(1.250000) ≈ 0.750000
			7'b0010101: sigmoid_out <= 7'b0001101;    //sigmoid(1.312500) ≈ 0.812500
			7'b0010110: sigmoid_out <= 7'b0001101;    //sigmoid(1.375000) ≈ 0.812500
			7'b0010111: sigmoid_out <= 7'b0001101;    //sigmoid(1.437500) ≈ 0.812500
			7'b0011000: sigmoid_out <= 7'b0001101;    //sigmoid(1.500000) ≈ 0.812500
			7'b0011001: sigmoid_out <= 7'b0001101;    //sigmoid(1.562500) ≈ 0.812500
			7'b0011010: sigmoid_out <= 7'b0001101;    //sigmoid(1.625000) ≈ 0.812500
			7'b0011011: sigmoid_out <= 7'b0001110;    //sigmoid(1.687500) ≈ 0.875000
			7'b0011100: sigmoid_out <= 7'b0001110;    //sigmoid(1.750000) ≈ 0.875000
			7'b0011101: sigmoid_out <= 7'b0001110;    //sigmoid(1.812500) ≈ 0.875000
			7'b0011110: sigmoid_out <= 7'b0001110;    //sigmoid(1.875000) ≈ 0.875000
			7'b0011111: sigmoid_out <= 7'b0001110;    //sigmoid(1.937500) ≈ 0.875000
			7'b0100000: sigmoid_out <= 7'b0001110;    //sigmoid(2.000000) ≈ 0.875000
			7'b0100001: sigmoid_out <= 7'b0001110;    //sigmoid(2.062500) ≈ 0.875000
			7'b0100010: sigmoid_out <= 7'b0001110;    //sigmoid(2.125000) ≈ 0.875000
			7'b0100011: sigmoid_out <= 7'b0001110;    //sigmoid(2.187500) ≈ 0.875000
			7'b0100100: sigmoid_out <= 7'b0001110;    //sigmoid(2.250000) ≈ 0.875000
			7'b0100101: sigmoid_out <= 7'b0001111;    //sigmoid(2.312500) ≈ 0.937500
			7'b0100110: sigmoid_out <= 7'b0001111;    //sigmoid(2.375000) ≈ 0.937500
			7'b0100111: sigmoid_out <= 7'b0001111;    //sigmoid(2.437500) ≈ 0.937500
			7'b0101000: sigmoid_out <= 7'b0001111;    //sigmoid(2.500000) ≈ 0.937500
			7'b0101001: sigmoid_out <= 7'b0001111;    //sigmoid(2.562500) ≈ 0.937500
			7'b0101010: sigmoid_out <= 7'b0001111;    //sigmoid(2.625000) ≈ 0.937500
			7'b0101011: sigmoid_out <= 7'b0001111;    //sigmoid(2.687500) ≈ 0.937500
			7'b0101100: sigmoid_out <= 7'b0001111;    //sigmoid(2.750000) ≈ 0.937500
			7'b0101101: sigmoid_out <= 7'b0001111;    //sigmoid(2.812500) ≈ 0.937500
			7'b0101110: sigmoid_out <= 7'b0001111;    //sigmoid(2.875000) ≈ 0.937500
			7'b0101111: sigmoid_out <= 7'b0001111;    //sigmoid(2.937500) ≈ 0.937500
			7'b0110000: sigmoid_out <= 7'b0001111;    //sigmoid(3.000000) ≈ 0.937500
			7'b0110001: sigmoid_out <= 7'b0001111;    //sigmoid(3.062500) ≈ 0.937500
			7'b0110010: sigmoid_out <= 7'b0001111;    //sigmoid(3.125000) ≈ 0.937500
			7'b0110011: sigmoid_out <= 7'b0001111;    //sigmoid(3.187500) ≈ 0.937500
			7'b0110100: sigmoid_out <= 7'b0001111;    //sigmoid(3.250000) ≈ 0.937500
			7'b0110101: sigmoid_out <= 7'b0001111;    //sigmoid(3.312500) ≈ 0.937500
			7'b0110110: sigmoid_out <= 7'b0001111;    //sigmoid(3.375000) ≈ 0.937500
			7'b0110111: sigmoid_out <= 7'b0010000;    //sigmoid(3.437500) ≈ 1.000000
			7'b0111000: sigmoid_out <= 7'b0010000;    //sigmoid(3.500000) ≈ 1.000000
			7'b0111001: sigmoid_out <= 7'b0010000;    //sigmoid(3.562500) ≈ 1.000000
			7'b0111010: sigmoid_out <= 7'b0010000;    //sigmoid(3.625000) ≈ 1.000000
			7'b0111011: sigmoid_out <= 7'b0010000;    //sigmoid(3.687500) ≈ 1.000000
			7'b0111100: sigmoid_out <= 7'b0010000;    //sigmoid(3.750000) ≈ 1.000000
			7'b0111101: sigmoid_out <= 7'b0010000;    //sigmoid(3.812500) ≈ 1.000000
			7'b0111110: sigmoid_out <= 7'b0010000;    //sigmoid(3.875000) ≈ 1.000000
			7'b0111111: sigmoid_out <= 7'b0010000;    //sigmoid(3.937500) ≈ 1.000000
			7'b1000000: sigmoid_out <= 7'b0010000;    //sigmoid(4.000000) ≈ 1.000000
			7'b1000001: sigmoid_out <= 7'b0010000;    //sigmoid(4.062500) ≈ 1.000000
			7'b1000010: sigmoid_out <= 7'b0010000;    //sigmoid(4.125000) ≈ 1.000000
			7'b1000011: sigmoid_out <= 7'b0010000;    //sigmoid(4.187500) ≈ 1.000000
			7'b1000100: sigmoid_out <= 7'b0010000;    //sigmoid(4.250000) ≈ 1.000000
			7'b1000101: sigmoid_out <= 7'b0010000;    //sigmoid(4.312500) ≈ 1.000000
			7'b1000110: sigmoid_out <= 7'b0010000;    //sigmoid(4.375000) ≈ 1.000000
			7'b1000111: sigmoid_out <= 7'b0010000;    //sigmoid(4.437500) ≈ 1.000000
			7'b1001000: sigmoid_out <= 7'b0010000;    //sigmoid(4.500000) ≈ 1.000000
			7'b1001001: sigmoid_out <= 7'b0010000;    //sigmoid(4.562500) ≈ 1.000000
			7'b1001010: sigmoid_out <= 7'b0010000;    //sigmoid(4.625000) ≈ 1.000000
			7'b1001011: sigmoid_out <= 7'b0010000;    //sigmoid(4.687500) ≈ 1.000000
			7'b1001100: sigmoid_out <= 7'b0010000;    //sigmoid(4.750000) ≈ 1.000000
			7'b1001101: sigmoid_out <= 7'b0010000;    //sigmoid(4.812500) ≈ 1.000000
			7'b1001110: sigmoid_out <= 7'b0010000;    //sigmoid(4.875000) ≈ 1.000000
			7'b1001111: sigmoid_out <= 7'b0010000;    //sigmoid(4.937500) ≈ 1.000000
			7'b1010000: sigmoid_out <= 7'b0010000;    //sigmoid(5.000000) ≈ 1.000000
			7'b1010001: sigmoid_out <= 7'b0010000;    //sigmoid(5.062500) ≈ 1.000000
			7'b1010010: sigmoid_out <= 7'b0010000;    //sigmoid(5.125000) ≈ 1.000000
			7'b1010011: sigmoid_out <= 7'b0010000;    //sigmoid(5.187500) ≈ 1.000000
			7'b1010100: sigmoid_out <= 7'b0010000;    //sigmoid(5.250000) ≈ 1.000000
			7'b1010101: sigmoid_out <= 7'b0010000;    //sigmoid(5.312500) ≈ 1.000000
			7'b1010110: sigmoid_out <= 7'b0010000;    //sigmoid(5.375000) ≈ 1.000000
			7'b1010111: sigmoid_out <= 7'b0010000;    //sigmoid(5.437500) ≈ 1.000000
			7'b1011000: sigmoid_out <= 7'b0010000;    //sigmoid(5.500000) ≈ 1.000000
			7'b1011001: sigmoid_out <= 7'b0010000;    //sigmoid(5.562500) ≈ 1.000000
			7'b1011010: sigmoid_out <= 7'b0010000;    //sigmoid(5.625000) ≈ 1.000000
			7'b1011011: sigmoid_out <= 7'b0010000;    //sigmoid(5.687500) ≈ 1.000000
			7'b1011100: sigmoid_out <= 7'b0010000;    //sigmoid(5.750000) ≈ 1.000000
			7'b1011101: sigmoid_out <= 7'b0010000;    //sigmoid(5.812500) ≈ 1.000000
			7'b1011110: sigmoid_out <= 7'b0010000;    //sigmoid(5.875000) ≈ 1.000000
			7'b1011111: sigmoid_out <= 7'b0010000;    //sigmoid(5.937500) ≈ 1.000000
			7'b1100000: sigmoid_out <= 7'b0010000;    //sigmoid(6.000000) ≈ 1.000000
			7'b1100001: sigmoid_out <= 7'b0010000;    //sigmoid(6.062500) ≈ 1.000000
			7'b1100010: sigmoid_out <= 7'b0010000;    //sigmoid(6.125000) ≈ 1.000000
			7'b1100011: sigmoid_out <= 7'b0010000;    //sigmoid(6.187500) ≈ 1.000000
			7'b1100100: sigmoid_out <= 7'b0010000;    //sigmoid(6.250000) ≈ 1.000000
			7'b1100101: sigmoid_out <= 7'b0010000;    //sigmoid(6.312500) ≈ 1.000000
			7'b1100110: sigmoid_out <= 7'b0010000;    //sigmoid(6.375000) ≈ 1.000000
			7'b1100111: sigmoid_out <= 7'b0010000;    //sigmoid(6.437500) ≈ 1.000000
			7'b1101000: sigmoid_out <= 7'b0010000;    //sigmoid(6.500000) ≈ 1.000000
			7'b1101001: sigmoid_out <= 7'b0010000;    //sigmoid(6.562500) ≈ 1.000000
			7'b1101010: sigmoid_out <= 7'b0010000;    //sigmoid(6.625000) ≈ 1.000000
			7'b1101011: sigmoid_out <= 7'b0010000;    //sigmoid(6.687500) ≈ 1.000000
			7'b1101100: sigmoid_out <= 7'b0010000;    //sigmoid(6.750000) ≈ 1.000000
			7'b1101101: sigmoid_out <= 7'b0010000;    //sigmoid(6.812500) ≈ 1.000000
			7'b1101110: sigmoid_out <= 7'b0010000;    //sigmoid(6.875000) ≈ 1.000000
			7'b1101111: sigmoid_out <= 7'b0010000;    //sigmoid(6.937500) ≈ 1.000000
			7'b1110000: sigmoid_out <= 7'b0010000;    //sigmoid(7.000000) ≈ 1.000000
			7'b1110001: sigmoid_out <= 7'b0010000;    //sigmoid(7.062500) ≈ 1.000000
			7'b1110010: sigmoid_out <= 7'b0010000;    //sigmoid(7.125000) ≈ 1.000000
			7'b1110011: sigmoid_out <= 7'b0010000;    //sigmoid(7.187500) ≈ 1.000000
			7'b1110100: sigmoid_out <= 7'b0010000;    //sigmoid(7.250000) ≈ 1.000000
			7'b1110101: sigmoid_out <= 7'b0010000;    //sigmoid(7.312500) ≈ 1.000000
			7'b1110110: sigmoid_out <= 7'b0010000;    //sigmoid(7.375000) ≈ 1.000000
			7'b1110111: sigmoid_out <= 7'b0010000;    //sigmoid(7.437500) ≈ 1.000000
			7'b1111000: sigmoid_out <= 7'b0010000;    //sigmoid(7.500000) ≈ 1.000000
			7'b1111001: sigmoid_out <= 7'b0010000;    //sigmoid(7.562500) ≈ 1.000000
			7'b1111010: sigmoid_out <= 7'b0010000;    //sigmoid(7.625000) ≈ 1.000000
			7'b1111011: sigmoid_out <= 7'b0010000;    //sigmoid(7.687500) ≈ 1.000000
			7'b1111100: sigmoid_out <= 7'b0010000;    //sigmoid(7.750000) ≈ 1.000000
			7'b1111101: sigmoid_out <= 7'b0010000;    //sigmoid(7.812500) ≈ 1.000000
			7'b1111110: sigmoid_out <= 7'b0010000;    //sigmoid(7.875000) ≈ 1.000000
			7'b1111111: sigmoid_out <= 7'b0010000;    //sigmoid(7.937500) ≈ 1.000000

        endcase
    end
endmodule