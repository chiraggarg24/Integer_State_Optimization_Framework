//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-06-28 14:36:01.428403
// Design Name: vanilla
// Module Name: sigmoidLUT_in7b3p_out9b8p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 7 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in7b3p_out9b8p #(
    parameter PRECISION_INPUT_BITS = 7,
    parameter PRECISION_OUTPUT_BITS = 9
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			7'b0000000: sigmoid_out <= 9'b010000000;    //sigmoid(0.000000) ≈ 0.500000
			7'b0000001: sigmoid_out <= 9'b010001000;    //sigmoid(0.125000) ≈ 0.531250
			7'b0000010: sigmoid_out <= 9'b010010000;    //sigmoid(0.250000) ≈ 0.562500
			7'b0000011: sigmoid_out <= 9'b010011000;    //sigmoid(0.375000) ≈ 0.593750
			7'b0000100: sigmoid_out <= 9'b010011111;    //sigmoid(0.500000) ≈ 0.621094
			7'b0000101: sigmoid_out <= 9'b010100111;    //sigmoid(0.625000) ≈ 0.652344
			7'b0000110: sigmoid_out <= 9'b010101110;    //sigmoid(0.750000) ≈ 0.679688
			7'b0000111: sigmoid_out <= 9'b010110101;    //sigmoid(0.875000) ≈ 0.707031
			7'b0001000: sigmoid_out <= 9'b010111011;    //sigmoid(1.000000) ≈ 0.730469
			7'b0001001: sigmoid_out <= 9'b011000001;    //sigmoid(1.125000) ≈ 0.753906
			7'b0001010: sigmoid_out <= 9'b011000111;    //sigmoid(1.250000) ≈ 0.777344
			7'b0001011: sigmoid_out <= 9'b011001100;    //sigmoid(1.375000) ≈ 0.796875
			7'b0001100: sigmoid_out <= 9'b011010001;    //sigmoid(1.500000) ≈ 0.816406
			7'b0001101: sigmoid_out <= 9'b011010110;    //sigmoid(1.625000) ≈ 0.835938
			7'b0001110: sigmoid_out <= 9'b011011010;    //sigmoid(1.750000) ≈ 0.851562
			7'b0001111: sigmoid_out <= 9'b011011110;    //sigmoid(1.875000) ≈ 0.867188
			7'b0010000: sigmoid_out <= 9'b011100001;    //sigmoid(2.000000) ≈ 0.878906
			7'b0010001: sigmoid_out <= 9'b011100101;    //sigmoid(2.125000) ≈ 0.894531
			7'b0010010: sigmoid_out <= 9'b011101000;    //sigmoid(2.250000) ≈ 0.906250
			7'b0010011: sigmoid_out <= 9'b011101010;    //sigmoid(2.375000) ≈ 0.914062
			7'b0010100: sigmoid_out <= 9'b011101101;    //sigmoid(2.500000) ≈ 0.925781
			7'b0010101: sigmoid_out <= 9'b011101111;    //sigmoid(2.625000) ≈ 0.933594
			7'b0010110: sigmoid_out <= 9'b011110001;    //sigmoid(2.750000) ≈ 0.941406
			7'b0010111: sigmoid_out <= 9'b011110010;    //sigmoid(2.875000) ≈ 0.945312
			7'b0011000: sigmoid_out <= 9'b011110100;    //sigmoid(3.000000) ≈ 0.953125
			7'b0011001: sigmoid_out <= 9'b011110101;    //sigmoid(3.125000) ≈ 0.957031
			7'b0011010: sigmoid_out <= 9'b011110110;    //sigmoid(3.250000) ≈ 0.960938
			7'b0011011: sigmoid_out <= 9'b011111000;    //sigmoid(3.375000) ≈ 0.968750
			7'b0011100: sigmoid_out <= 9'b011111000;    //sigmoid(3.500000) ≈ 0.968750
			7'b0011101: sigmoid_out <= 9'b011111001;    //sigmoid(3.625000) ≈ 0.972656
			7'b0011110: sigmoid_out <= 9'b011111010;    //sigmoid(3.750000) ≈ 0.976562
			7'b0011111: sigmoid_out <= 9'b011111011;    //sigmoid(3.875000) ≈ 0.980469
			7'b0100000: sigmoid_out <= 9'b011111011;    //sigmoid(4.000000) ≈ 0.980469
			7'b0100001: sigmoid_out <= 9'b011111100;    //sigmoid(4.125000) ≈ 0.984375
			7'b0100010: sigmoid_out <= 9'b011111100;    //sigmoid(4.250000) ≈ 0.984375
			7'b0100011: sigmoid_out <= 9'b011111101;    //sigmoid(4.375000) ≈ 0.988281
			7'b0100100: sigmoid_out <= 9'b011111101;    //sigmoid(4.500000) ≈ 0.988281
			7'b0100101: sigmoid_out <= 9'b011111110;    //sigmoid(4.625000) ≈ 0.992188
			7'b0100110: sigmoid_out <= 9'b011111110;    //sigmoid(4.750000) ≈ 0.992188
			7'b0100111: sigmoid_out <= 9'b011111110;    //sigmoid(4.875000) ≈ 0.992188
			7'b0101000: sigmoid_out <= 9'b011111110;    //sigmoid(5.000000) ≈ 0.992188
			7'b0101001: sigmoid_out <= 9'b011111110;    //sigmoid(5.125000) ≈ 0.992188
			7'b0101010: sigmoid_out <= 9'b011111111;    //sigmoid(5.250000) ≈ 0.996094
			7'b0101011: sigmoid_out <= 9'b011111111;    //sigmoid(5.375000) ≈ 0.996094
			7'b0101100: sigmoid_out <= 9'b011111111;    //sigmoid(5.500000) ≈ 0.996094
			7'b0101101: sigmoid_out <= 9'b011111111;    //sigmoid(5.625000) ≈ 0.996094
			7'b0101110: sigmoid_out <= 9'b011111111;    //sigmoid(5.750000) ≈ 0.996094
			7'b0101111: sigmoid_out <= 9'b011111111;    //sigmoid(5.875000) ≈ 0.996094
			7'b0110000: sigmoid_out <= 9'b011111111;    //sigmoid(6.000000) ≈ 0.996094
			7'b0110001: sigmoid_out <= 9'b011111111;    //sigmoid(6.125000) ≈ 0.996094
			7'b0110010: sigmoid_out <= 9'b100000000;    //sigmoid(6.250000) ≈ 1.000000
			7'b0110011: sigmoid_out <= 9'b100000000;    //sigmoid(6.375000) ≈ 1.000000
			7'b0110100: sigmoid_out <= 9'b100000000;    //sigmoid(6.500000) ≈ 1.000000
			7'b0110101: sigmoid_out <= 9'b100000000;    //sigmoid(6.625000) ≈ 1.000000
			7'b0110110: sigmoid_out <= 9'b100000000;    //sigmoid(6.750000) ≈ 1.000000
			7'b0110111: sigmoid_out <= 9'b100000000;    //sigmoid(6.875000) ≈ 1.000000
			7'b0111000: sigmoid_out <= 9'b100000000;    //sigmoid(7.000000) ≈ 1.000000
			7'b0111001: sigmoid_out <= 9'b100000000;    //sigmoid(7.125000) ≈ 1.000000
			7'b0111010: sigmoid_out <= 9'b100000000;    //sigmoid(7.250000) ≈ 1.000000
			7'b0111011: sigmoid_out <= 9'b100000000;    //sigmoid(7.375000) ≈ 1.000000
			7'b0111100: sigmoid_out <= 9'b100000000;    //sigmoid(7.500000) ≈ 1.000000
			7'b0111101: sigmoid_out <= 9'b100000000;    //sigmoid(7.625000) ≈ 1.000000
			7'b0111110: sigmoid_out <= 9'b100000000;    //sigmoid(7.750000) ≈ 1.000000
			7'b0111111: sigmoid_out <= 9'b100000000;    //sigmoid(7.875000) ≈ 1.000000
			7'b1000000: sigmoid_out <= 9'b100000000;    //sigmoid(8.000000) ≈ 1.000000
			7'b1000001: sigmoid_out <= 9'b100000000;    //sigmoid(8.125000) ≈ 1.000000
			7'b1000010: sigmoid_out <= 9'b100000000;    //sigmoid(8.250000) ≈ 1.000000
			7'b1000011: sigmoid_out <= 9'b100000000;    //sigmoid(8.375000) ≈ 1.000000
			7'b1000100: sigmoid_out <= 9'b100000000;    //sigmoid(8.500000) ≈ 1.000000
			7'b1000101: sigmoid_out <= 9'b100000000;    //sigmoid(8.625000) ≈ 1.000000
			7'b1000110: sigmoid_out <= 9'b100000000;    //sigmoid(8.750000) ≈ 1.000000
			7'b1000111: sigmoid_out <= 9'b100000000;    //sigmoid(8.875000) ≈ 1.000000
			7'b1001000: sigmoid_out <= 9'b100000000;    //sigmoid(9.000000) ≈ 1.000000
			7'b1001001: sigmoid_out <= 9'b100000000;    //sigmoid(9.125000) ≈ 1.000000
			7'b1001010: sigmoid_out <= 9'b100000000;    //sigmoid(9.250000) ≈ 1.000000
			7'b1001011: sigmoid_out <= 9'b100000000;    //sigmoid(9.375000) ≈ 1.000000
			7'b1001100: sigmoid_out <= 9'b100000000;    //sigmoid(9.500000) ≈ 1.000000
			7'b1001101: sigmoid_out <= 9'b100000000;    //sigmoid(9.625000) ≈ 1.000000
			7'b1001110: sigmoid_out <= 9'b100000000;    //sigmoid(9.750000) ≈ 1.000000
			7'b1001111: sigmoid_out <= 9'b100000000;    //sigmoid(9.875000) ≈ 1.000000
			7'b1010000: sigmoid_out <= 9'b100000000;    //sigmoid(10.000000) ≈ 1.000000
			7'b1010001: sigmoid_out <= 9'b100000000;    //sigmoid(10.125000) ≈ 1.000000
			7'b1010010: sigmoid_out <= 9'b100000000;    //sigmoid(10.250000) ≈ 1.000000
			7'b1010011: sigmoid_out <= 9'b100000000;    //sigmoid(10.375000) ≈ 1.000000
			7'b1010100: sigmoid_out <= 9'b100000000;    //sigmoid(10.500000) ≈ 1.000000
			7'b1010101: sigmoid_out <= 9'b100000000;    //sigmoid(10.625000) ≈ 1.000000
			7'b1010110: sigmoid_out <= 9'b100000000;    //sigmoid(10.750000) ≈ 1.000000
			7'b1010111: sigmoid_out <= 9'b100000000;    //sigmoid(10.875000) ≈ 1.000000
			7'b1011000: sigmoid_out <= 9'b100000000;    //sigmoid(11.000000) ≈ 1.000000
			7'b1011001: sigmoid_out <= 9'b100000000;    //sigmoid(11.125000) ≈ 1.000000
			7'b1011010: sigmoid_out <= 9'b100000000;    //sigmoid(11.250000) ≈ 1.000000
			7'b1011011: sigmoid_out <= 9'b100000000;    //sigmoid(11.375000) ≈ 1.000000
			7'b1011100: sigmoid_out <= 9'b100000000;    //sigmoid(11.500000) ≈ 1.000000
			7'b1011101: sigmoid_out <= 9'b100000000;    //sigmoid(11.625000) ≈ 1.000000
			7'b1011110: sigmoid_out <= 9'b100000000;    //sigmoid(11.750000) ≈ 1.000000
			7'b1011111: sigmoid_out <= 9'b100000000;    //sigmoid(11.875000) ≈ 1.000000
			7'b1100000: sigmoid_out <= 9'b100000000;    //sigmoid(12.000000) ≈ 1.000000
			7'b1100001: sigmoid_out <= 9'b100000000;    //sigmoid(12.125000) ≈ 1.000000
			7'b1100010: sigmoid_out <= 9'b100000000;    //sigmoid(12.250000) ≈ 1.000000
			7'b1100011: sigmoid_out <= 9'b100000000;    //sigmoid(12.375000) ≈ 1.000000
			7'b1100100: sigmoid_out <= 9'b100000000;    //sigmoid(12.500000) ≈ 1.000000
			7'b1100101: sigmoid_out <= 9'b100000000;    //sigmoid(12.625000) ≈ 1.000000
			7'b1100110: sigmoid_out <= 9'b100000000;    //sigmoid(12.750000) ≈ 1.000000
			7'b1100111: sigmoid_out <= 9'b100000000;    //sigmoid(12.875000) ≈ 1.000000
			7'b1101000: sigmoid_out <= 9'b100000000;    //sigmoid(13.000000) ≈ 1.000000
			7'b1101001: sigmoid_out <= 9'b100000000;    //sigmoid(13.125000) ≈ 1.000000
			7'b1101010: sigmoid_out <= 9'b100000000;    //sigmoid(13.250000) ≈ 1.000000
			7'b1101011: sigmoid_out <= 9'b100000000;    //sigmoid(13.375000) ≈ 1.000000
			7'b1101100: sigmoid_out <= 9'b100000000;    //sigmoid(13.500000) ≈ 1.000000
			7'b1101101: sigmoid_out <= 9'b100000000;    //sigmoid(13.625000) ≈ 1.000000
			7'b1101110: sigmoid_out <= 9'b100000000;    //sigmoid(13.750000) ≈ 1.000000
			7'b1101111: sigmoid_out <= 9'b100000000;    //sigmoid(13.875000) ≈ 1.000000
			7'b1110000: sigmoid_out <= 9'b100000000;    //sigmoid(14.000000) ≈ 1.000000
			7'b1110001: sigmoid_out <= 9'b100000000;    //sigmoid(14.125000) ≈ 1.000000
			7'b1110010: sigmoid_out <= 9'b100000000;    //sigmoid(14.250000) ≈ 1.000000
			7'b1110011: sigmoid_out <= 9'b100000000;    //sigmoid(14.375000) ≈ 1.000000
			7'b1110100: sigmoid_out <= 9'b100000000;    //sigmoid(14.500000) ≈ 1.000000
			7'b1110101: sigmoid_out <= 9'b100000000;    //sigmoid(14.625000) ≈ 1.000000
			7'b1110110: sigmoid_out <= 9'b100000000;    //sigmoid(14.750000) ≈ 1.000000
			7'b1110111: sigmoid_out <= 9'b100000000;    //sigmoid(14.875000) ≈ 1.000000
			7'b1111000: sigmoid_out <= 9'b100000000;    //sigmoid(15.000000) ≈ 1.000000
			7'b1111001: sigmoid_out <= 9'b100000000;    //sigmoid(15.125000) ≈ 1.000000
			7'b1111010: sigmoid_out <= 9'b100000000;    //sigmoid(15.250000) ≈ 1.000000
			7'b1111011: sigmoid_out <= 9'b100000000;    //sigmoid(15.375000) ≈ 1.000000
			7'b1111100: sigmoid_out <= 9'b100000000;    //sigmoid(15.500000) ≈ 1.000000
			7'b1111101: sigmoid_out <= 9'b100000000;    //sigmoid(15.625000) ≈ 1.000000
			7'b1111110: sigmoid_out <= 9'b100000000;    //sigmoid(15.750000) ≈ 1.000000
			7'b1111111: sigmoid_out <= 9'b100000000;    //sigmoid(15.875000) ≈ 1.000000

        endcase
    end
endmodule