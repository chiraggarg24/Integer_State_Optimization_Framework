//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
//
// Create Date: 2019-06-28 15:31:06.522243
// Design Name: vanilla
// Module Name: sigmoidLUT_in7b4p_out12b11p
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 7 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
//
// Additional Comments: Generated by LUT_generator_sigmoid.py
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_in7b4p_out12b11p #(
    parameter PRECISION_INPUT_BITS = 7,
    parameter PRECISION_OUTPUT_BITS = 12
)(
    input[PRECISION_INPUT_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_OUTPUT_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			7'b0000000: sigmoid_out <= 12'b010000000000;    //sigmoid(0.000000) ≈ 0.500000
			7'b0000001: sigmoid_out <= 12'b010000100000;    //sigmoid(0.062500) ≈ 0.515625
			7'b0000010: sigmoid_out <= 12'b010001000000;    //sigmoid(0.125000) ≈ 0.531250
			7'b0000011: sigmoid_out <= 12'b010001100000;    //sigmoid(0.187500) ≈ 0.546875
			7'b0000100: sigmoid_out <= 12'b010001111111;    //sigmoid(0.250000) ≈ 0.562012
			7'b0000101: sigmoid_out <= 12'b010010011111;    //sigmoid(0.312500) ≈ 0.577637
			7'b0000110: sigmoid_out <= 12'b010010111110;    //sigmoid(0.375000) ≈ 0.592773
			7'b0000111: sigmoid_out <= 12'b010011011100;    //sigmoid(0.437500) ≈ 0.607422
			7'b0001000: sigmoid_out <= 12'b010011111011;    //sigmoid(0.500000) ≈ 0.622559
			7'b0001001: sigmoid_out <= 12'b010100011001;    //sigmoid(0.562500) ≈ 0.637207
			7'b0001010: sigmoid_out <= 12'b010100110110;    //sigmoid(0.625000) ≈ 0.651367
			7'b0001011: sigmoid_out <= 12'b010101010011;    //sigmoid(0.687500) ≈ 0.665527
			7'b0001100: sigmoid_out <= 12'b010101101111;    //sigmoid(0.750000) ≈ 0.679199
			7'b0001101: sigmoid_out <= 12'b010110001011;    //sigmoid(0.812500) ≈ 0.692871
			7'b0001110: sigmoid_out <= 12'b010110100101;    //sigmoid(0.875000) ≈ 0.705566
			7'b0001111: sigmoid_out <= 12'b010111000000;    //sigmoid(0.937500) ≈ 0.718750
			7'b0010000: sigmoid_out <= 12'b010111011001;    //sigmoid(1.000000) ≈ 0.730957
			7'b0010001: sigmoid_out <= 12'b010111110010;    //sigmoid(1.062500) ≈ 0.743164
			7'b0010010: sigmoid_out <= 12'b011000001010;    //sigmoid(1.125000) ≈ 0.754883
			7'b0010011: sigmoid_out <= 12'b011000100001;    //sigmoid(1.187500) ≈ 0.766113
			7'b0010100: sigmoid_out <= 12'b011000111000;    //sigmoid(1.250000) ≈ 0.777344
			7'b0010101: sigmoid_out <= 12'b011001001110;    //sigmoid(1.312500) ≈ 0.788086
			7'b0010110: sigmoid_out <= 12'b011001100011;    //sigmoid(1.375000) ≈ 0.798340
			7'b0010111: sigmoid_out <= 12'b011001110111;    //sigmoid(1.437500) ≈ 0.808105
			7'b0011000: sigmoid_out <= 12'b011010001010;    //sigmoid(1.500000) ≈ 0.817383
			7'b0011001: sigmoid_out <= 12'b011010011101;    //sigmoid(1.562500) ≈ 0.826660
			7'b0011010: sigmoid_out <= 12'b011010101111;    //sigmoid(1.625000) ≈ 0.835449
			7'b0011011: sigmoid_out <= 12'b011011000000;    //sigmoid(1.687500) ≈ 0.843750
			7'b0011100: sigmoid_out <= 12'b011011010001;    //sigmoid(1.750000) ≈ 0.852051
			7'b0011101: sigmoid_out <= 12'b011011100001;    //sigmoid(1.812500) ≈ 0.859863
			7'b0011110: sigmoid_out <= 12'b011011110000;    //sigmoid(1.875000) ≈ 0.867188
			7'b0011111: sigmoid_out <= 12'b011011111110;    //sigmoid(1.937500) ≈ 0.874023
			7'b0100000: sigmoid_out <= 12'b011100001100;    //sigmoid(2.000000) ≈ 0.880859
			7'b0100001: sigmoid_out <= 12'b011100011001;    //sigmoid(2.062500) ≈ 0.887207
			7'b0100010: sigmoid_out <= 12'b011100100101;    //sigmoid(2.125000) ≈ 0.893066
			7'b0100011: sigmoid_out <= 12'b011100110001;    //sigmoid(2.187500) ≈ 0.898926
			7'b0100100: sigmoid_out <= 12'b011100111101;    //sigmoid(2.250000) ≈ 0.904785
			7'b0100101: sigmoid_out <= 12'b011101000111;    //sigmoid(2.312500) ≈ 0.909668
			7'b0100110: sigmoid_out <= 12'b011101010010;    //sigmoid(2.375000) ≈ 0.915039
			7'b0100111: sigmoid_out <= 12'b011101011011;    //sigmoid(2.437500) ≈ 0.919434
			7'b0101000: sigmoid_out <= 12'b011101100101;    //sigmoid(2.500000) ≈ 0.924316
			7'b0101001: sigmoid_out <= 12'b011101101101;    //sigmoid(2.562500) ≈ 0.928223
			7'b0101010: sigmoid_out <= 12'b011101110110;    //sigmoid(2.625000) ≈ 0.932617
			7'b0101011: sigmoid_out <= 12'b011101111110;    //sigmoid(2.687500) ≈ 0.936523
			7'b0101100: sigmoid_out <= 12'b011110000101;    //sigmoid(2.750000) ≈ 0.939941
			7'b0101101: sigmoid_out <= 12'b011110001100;    //sigmoid(2.812500) ≈ 0.943359
			7'b0101110: sigmoid_out <= 12'b011110010011;    //sigmoid(2.875000) ≈ 0.946777
			7'b0101111: sigmoid_out <= 12'b011110011001;    //sigmoid(2.937500) ≈ 0.949707
			7'b0110000: sigmoid_out <= 12'b011110011111;    //sigmoid(3.000000) ≈ 0.952637
			7'b0110001: sigmoid_out <= 12'b011110100100;    //sigmoid(3.062500) ≈ 0.955078
			7'b0110010: sigmoid_out <= 12'b011110101010;    //sigmoid(3.125000) ≈ 0.958008
			7'b0110011: sigmoid_out <= 12'b011110101111;    //sigmoid(3.187500) ≈ 0.960449
			7'b0110100: sigmoid_out <= 12'b011110110100;    //sigmoid(3.250000) ≈ 0.962891
			7'b0110101: sigmoid_out <= 12'b011110111000;    //sigmoid(3.312500) ≈ 0.964844
			7'b0110110: sigmoid_out <= 12'b011110111100;    //sigmoid(3.375000) ≈ 0.966797
			7'b0110111: sigmoid_out <= 12'b011111000000;    //sigmoid(3.437500) ≈ 0.968750
			7'b0111000: sigmoid_out <= 12'b011111000100;    //sigmoid(3.500000) ≈ 0.970703
			7'b0111001: sigmoid_out <= 12'b011111001000;    //sigmoid(3.562500) ≈ 0.972656
			7'b0111010: sigmoid_out <= 12'b011111001011;    //sigmoid(3.625000) ≈ 0.974121
			7'b0111011: sigmoid_out <= 12'b011111001110;    //sigmoid(3.687500) ≈ 0.975586
			7'b0111100: sigmoid_out <= 12'b011111010001;    //sigmoid(3.750000) ≈ 0.977051
			7'b0111101: sigmoid_out <= 12'b011111010100;    //sigmoid(3.812500) ≈ 0.978516
			7'b0111110: sigmoid_out <= 12'b011111010110;    //sigmoid(3.875000) ≈ 0.979492
			7'b0111111: sigmoid_out <= 12'b011111011001;    //sigmoid(3.937500) ≈ 0.980957
			7'b1000000: sigmoid_out <= 12'b011111011011;    //sigmoid(4.000000) ≈ 0.981934
			7'b1000001: sigmoid_out <= 12'b011111011101;    //sigmoid(4.062500) ≈ 0.982910
			7'b1000010: sigmoid_out <= 12'b011111011111;    //sigmoid(4.125000) ≈ 0.983887
			7'b1000011: sigmoid_out <= 12'b011111100001;    //sigmoid(4.187500) ≈ 0.984863
			7'b1000100: sigmoid_out <= 12'b011111100011;    //sigmoid(4.250000) ≈ 0.985840
			7'b1000101: sigmoid_out <= 12'b011111100101;    //sigmoid(4.312500) ≈ 0.986816
			7'b1000110: sigmoid_out <= 12'b011111100111;    //sigmoid(4.375000) ≈ 0.987793
			7'b1000111: sigmoid_out <= 12'b011111101000;    //sigmoid(4.437500) ≈ 0.988281
			7'b1001000: sigmoid_out <= 12'b011111101001;    //sigmoid(4.500000) ≈ 0.988770
			7'b1001001: sigmoid_out <= 12'b011111101011;    //sigmoid(4.562500) ≈ 0.989746
			7'b1001010: sigmoid_out <= 12'b011111101100;    //sigmoid(4.625000) ≈ 0.990234
			7'b1001011: sigmoid_out <= 12'b011111101101;    //sigmoid(4.687500) ≈ 0.990723
			7'b1001100: sigmoid_out <= 12'b011111101110;    //sigmoid(4.750000) ≈ 0.991211
			7'b1001101: sigmoid_out <= 12'b011111101111;    //sigmoid(4.812500) ≈ 0.991699
			7'b1001110: sigmoid_out <= 12'b011111110000;    //sigmoid(4.875000) ≈ 0.992188
			7'b1001111: sigmoid_out <= 12'b011111110001;    //sigmoid(4.937500) ≈ 0.992676
			7'b1010000: sigmoid_out <= 12'b011111110010;    //sigmoid(5.000000) ≈ 0.993164
			7'b1010001: sigmoid_out <= 12'b011111110011;    //sigmoid(5.062500) ≈ 0.993652
			7'b1010010: sigmoid_out <= 12'b011111110100;    //sigmoid(5.125000) ≈ 0.994141
			7'b1010011: sigmoid_out <= 12'b011111110101;    //sigmoid(5.187500) ≈ 0.994629
			7'b1010100: sigmoid_out <= 12'b011111110101;    //sigmoid(5.250000) ≈ 0.994629
			7'b1010101: sigmoid_out <= 12'b011111110110;    //sigmoid(5.312500) ≈ 0.995117
			7'b1010110: sigmoid_out <= 12'b011111110111;    //sigmoid(5.375000) ≈ 0.995605
			7'b1010111: sigmoid_out <= 12'b011111110111;    //sigmoid(5.437500) ≈ 0.995605
			7'b1011000: sigmoid_out <= 12'b011111111000;    //sigmoid(5.500000) ≈ 0.996094
			7'b1011001: sigmoid_out <= 12'b011111111000;    //sigmoid(5.562500) ≈ 0.996094
			7'b1011010: sigmoid_out <= 12'b011111111001;    //sigmoid(5.625000) ≈ 0.996582
			7'b1011011: sigmoid_out <= 12'b011111111001;    //sigmoid(5.687500) ≈ 0.996582
			7'b1011100: sigmoid_out <= 12'b011111111010;    //sigmoid(5.750000) ≈ 0.997070
			7'b1011101: sigmoid_out <= 12'b011111111010;    //sigmoid(5.812500) ≈ 0.997070
			7'b1011110: sigmoid_out <= 12'b011111111010;    //sigmoid(5.875000) ≈ 0.997070
			7'b1011111: sigmoid_out <= 12'b011111111011;    //sigmoid(5.937500) ≈ 0.997559
			7'b1100000: sigmoid_out <= 12'b011111111011;    //sigmoid(6.000000) ≈ 0.997559
			7'b1100001: sigmoid_out <= 12'b011111111011;    //sigmoid(6.062500) ≈ 0.997559
			7'b1100010: sigmoid_out <= 12'b011111111100;    //sigmoid(6.125000) ≈ 0.998047
			7'b1100011: sigmoid_out <= 12'b011111111100;    //sigmoid(6.187500) ≈ 0.998047
			7'b1100100: sigmoid_out <= 12'b011111111100;    //sigmoid(6.250000) ≈ 0.998047
			7'b1100101: sigmoid_out <= 12'b011111111100;    //sigmoid(6.312500) ≈ 0.998047
			7'b1100110: sigmoid_out <= 12'b011111111101;    //sigmoid(6.375000) ≈ 0.998535
			7'b1100111: sigmoid_out <= 12'b011111111101;    //sigmoid(6.437500) ≈ 0.998535
			7'b1101000: sigmoid_out <= 12'b011111111101;    //sigmoid(6.500000) ≈ 0.998535
			7'b1101001: sigmoid_out <= 12'b011111111101;    //sigmoid(6.562500) ≈ 0.998535
			7'b1101010: sigmoid_out <= 12'b011111111101;    //sigmoid(6.625000) ≈ 0.998535
			7'b1101011: sigmoid_out <= 12'b011111111101;    //sigmoid(6.687500) ≈ 0.998535
			7'b1101100: sigmoid_out <= 12'b011111111110;    //sigmoid(6.750000) ≈ 0.999023
			7'b1101101: sigmoid_out <= 12'b011111111110;    //sigmoid(6.812500) ≈ 0.999023
			7'b1101110: sigmoid_out <= 12'b011111111110;    //sigmoid(6.875000) ≈ 0.999023
			7'b1101111: sigmoid_out <= 12'b011111111110;    //sigmoid(6.937500) ≈ 0.999023
			7'b1110000: sigmoid_out <= 12'b011111111110;    //sigmoid(7.000000) ≈ 0.999023
			7'b1110001: sigmoid_out <= 12'b011111111110;    //sigmoid(7.062500) ≈ 0.999023
			7'b1110010: sigmoid_out <= 12'b011111111110;    //sigmoid(7.125000) ≈ 0.999023
			7'b1110011: sigmoid_out <= 12'b011111111110;    //sigmoid(7.187500) ≈ 0.999023
			7'b1110100: sigmoid_out <= 12'b011111111111;    //sigmoid(7.250000) ≈ 0.999512
			7'b1110101: sigmoid_out <= 12'b011111111111;    //sigmoid(7.312500) ≈ 0.999512
			7'b1110110: sigmoid_out <= 12'b011111111111;    //sigmoid(7.375000) ≈ 0.999512
			7'b1110111: sigmoid_out <= 12'b011111111111;    //sigmoid(7.437500) ≈ 0.999512
			7'b1111000: sigmoid_out <= 12'b011111111111;    //sigmoid(7.500000) ≈ 0.999512
			7'b1111001: sigmoid_out <= 12'b011111111111;    //sigmoid(7.562500) ≈ 0.999512
			7'b1111010: sigmoid_out <= 12'b011111111111;    //sigmoid(7.625000) ≈ 0.999512
			7'b1111011: sigmoid_out <= 12'b011111111111;    //sigmoid(7.687500) ≈ 0.999512
			7'b1111100: sigmoid_out <= 12'b011111111111;    //sigmoid(7.750000) ≈ 0.999512
			7'b1111101: sigmoid_out <= 12'b011111111111;    //sigmoid(7.812500) ≈ 0.999512
			7'b1111110: sigmoid_out <= 12'b011111111111;    //sigmoid(7.875000) ≈ 0.999512
			7'b1111111: sigmoid_out <= 12'b011111111111;    //sigmoid(7.937500) ≈ 0.999512

        endcase
    end
endmodule