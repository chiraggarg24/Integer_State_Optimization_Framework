//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
// 
// Create Date: 2019-06-28 14:19:00.068336
// Design Name: vanilla
// Module Name: sigmoidLUT_9bit_5point
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 9 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
// 
// Additional Comments: Generated by LUT_generator_sigmoid.py
// 
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_9bit_5point #(
    parameter PRECISION_BITS = 9
)(
    input[PRECISION_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			9'b000000000: sigmoid_out <= 9'b000010000;    //sigmoid(0.000000) ≈ 0.500000
			9'b000000001: sigmoid_out <= 9'b000010000;    //sigmoid(0.031250) ≈ 0.500000
			9'b000000010: sigmoid_out <= 9'b000010000;    //sigmoid(0.062500) ≈ 0.500000
			9'b000000011: sigmoid_out <= 9'b000010001;    //sigmoid(0.093750) ≈ 0.531250
			9'b000000100: sigmoid_out <= 9'b000010001;    //sigmoid(0.125000) ≈ 0.531250
			9'b000000101: sigmoid_out <= 9'b000010001;    //sigmoid(0.156250) ≈ 0.531250
			9'b000000110: sigmoid_out <= 9'b000010001;    //sigmoid(0.187500) ≈ 0.531250
			9'b000000111: sigmoid_out <= 9'b000010010;    //sigmoid(0.218750) ≈ 0.562500
			9'b000001000: sigmoid_out <= 9'b000010010;    //sigmoid(0.250000) ≈ 0.562500
			9'b000001001: sigmoid_out <= 9'b000010010;    //sigmoid(0.281250) ≈ 0.562500
			9'b000001010: sigmoid_out <= 9'b000010010;    //sigmoid(0.312500) ≈ 0.562500
			9'b000001011: sigmoid_out <= 9'b000010011;    //sigmoid(0.343750) ≈ 0.593750
			9'b000001100: sigmoid_out <= 9'b000010011;    //sigmoid(0.375000) ≈ 0.593750
			9'b000001101: sigmoid_out <= 9'b000010011;    //sigmoid(0.406250) ≈ 0.593750
			9'b000001110: sigmoid_out <= 9'b000010011;    //sigmoid(0.437500) ≈ 0.593750
			9'b000001111: sigmoid_out <= 9'b000010100;    //sigmoid(0.468750) ≈ 0.625000
			9'b000010000: sigmoid_out <= 9'b000010100;    //sigmoid(0.500000) ≈ 0.625000
			9'b000010001: sigmoid_out <= 9'b000010100;    //sigmoid(0.531250) ≈ 0.625000
			9'b000010010: sigmoid_out <= 9'b000010100;    //sigmoid(0.562500) ≈ 0.625000
			9'b000010011: sigmoid_out <= 9'b000010101;    //sigmoid(0.593750) ≈ 0.656250
			9'b000010100: sigmoid_out <= 9'b000010101;    //sigmoid(0.625000) ≈ 0.656250
			9'b000010101: sigmoid_out <= 9'b000010101;    //sigmoid(0.656250) ≈ 0.656250
			9'b000010110: sigmoid_out <= 9'b000010101;    //sigmoid(0.687500) ≈ 0.656250
			9'b000010111: sigmoid_out <= 9'b000010110;    //sigmoid(0.718750) ≈ 0.687500
			9'b000011000: sigmoid_out <= 9'b000010110;    //sigmoid(0.750000) ≈ 0.687500
			9'b000011001: sigmoid_out <= 9'b000010110;    //sigmoid(0.781250) ≈ 0.687500
			9'b000011010: sigmoid_out <= 9'b000010110;    //sigmoid(0.812500) ≈ 0.687500
			9'b000011011: sigmoid_out <= 9'b000010110;    //sigmoid(0.843750) ≈ 0.687500
			9'b000011100: sigmoid_out <= 9'b000010111;    //sigmoid(0.875000) ≈ 0.718750
			9'b000011101: sigmoid_out <= 9'b000010111;    //sigmoid(0.906250) ≈ 0.718750
			9'b000011110: sigmoid_out <= 9'b000010111;    //sigmoid(0.937500) ≈ 0.718750
			9'b000011111: sigmoid_out <= 9'b000010111;    //sigmoid(0.968750) ≈ 0.718750
			9'b000100000: sigmoid_out <= 9'b000010111;    //sigmoid(1.000000) ≈ 0.718750
			9'b000100001: sigmoid_out <= 9'b000011000;    //sigmoid(1.031250) ≈ 0.750000
			9'b000100010: sigmoid_out <= 9'b000011000;    //sigmoid(1.062500) ≈ 0.750000
			9'b000100011: sigmoid_out <= 9'b000011000;    //sigmoid(1.093750) ≈ 0.750000
			9'b000100100: sigmoid_out <= 9'b000011000;    //sigmoid(1.125000) ≈ 0.750000
			9'b000100101: sigmoid_out <= 9'b000011000;    //sigmoid(1.156250) ≈ 0.750000
			9'b000100110: sigmoid_out <= 9'b000011001;    //sigmoid(1.187500) ≈ 0.781250
			9'b000100111: sigmoid_out <= 9'b000011001;    //sigmoid(1.218750) ≈ 0.781250
			9'b000101000: sigmoid_out <= 9'b000011001;    //sigmoid(1.250000) ≈ 0.781250
			9'b000101001: sigmoid_out <= 9'b000011001;    //sigmoid(1.281250) ≈ 0.781250
			9'b000101010: sigmoid_out <= 9'b000011001;    //sigmoid(1.312500) ≈ 0.781250
			9'b000101011: sigmoid_out <= 9'b000011001;    //sigmoid(1.343750) ≈ 0.781250
			9'b000101100: sigmoid_out <= 9'b000011010;    //sigmoid(1.375000) ≈ 0.812500
			9'b000101101: sigmoid_out <= 9'b000011010;    //sigmoid(1.406250) ≈ 0.812500
			9'b000101110: sigmoid_out <= 9'b000011010;    //sigmoid(1.437500) ≈ 0.812500
			9'b000101111: sigmoid_out <= 9'b000011010;    //sigmoid(1.468750) ≈ 0.812500
			9'b000110000: sigmoid_out <= 9'b000011010;    //sigmoid(1.500000) ≈ 0.812500
			9'b000110001: sigmoid_out <= 9'b000011010;    //sigmoid(1.531250) ≈ 0.812500
			9'b000110010: sigmoid_out <= 9'b000011010;    //sigmoid(1.562500) ≈ 0.812500
			9'b000110011: sigmoid_out <= 9'b000011011;    //sigmoid(1.593750) ≈ 0.843750
			9'b000110100: sigmoid_out <= 9'b000011011;    //sigmoid(1.625000) ≈ 0.843750
			9'b000110101: sigmoid_out <= 9'b000011011;    //sigmoid(1.656250) ≈ 0.843750
			9'b000110110: sigmoid_out <= 9'b000011011;    //sigmoid(1.687500) ≈ 0.843750
			9'b000110111: sigmoid_out <= 9'b000011011;    //sigmoid(1.718750) ≈ 0.843750
			9'b000111000: sigmoid_out <= 9'b000011011;    //sigmoid(1.750000) ≈ 0.843750
			9'b000111001: sigmoid_out <= 9'b000011011;    //sigmoid(1.781250) ≈ 0.843750
			9'b000111010: sigmoid_out <= 9'b000011100;    //sigmoid(1.812500) ≈ 0.875000
			9'b000111011: sigmoid_out <= 9'b000011100;    //sigmoid(1.843750) ≈ 0.875000
			9'b000111100: sigmoid_out <= 9'b000011100;    //sigmoid(1.875000) ≈ 0.875000
			9'b000111101: sigmoid_out <= 9'b000011100;    //sigmoid(1.906250) ≈ 0.875000
			9'b000111110: sigmoid_out <= 9'b000011100;    //sigmoid(1.937500) ≈ 0.875000
			9'b000111111: sigmoid_out <= 9'b000011100;    //sigmoid(1.968750) ≈ 0.875000
			9'b001000000: sigmoid_out <= 9'b000011100;    //sigmoid(2.000000) ≈ 0.875000
			9'b001000001: sigmoid_out <= 9'b000011100;    //sigmoid(2.031250) ≈ 0.875000
			9'b001000010: sigmoid_out <= 9'b000011100;    //sigmoid(2.062500) ≈ 0.875000
			9'b001000011: sigmoid_out <= 9'b000011100;    //sigmoid(2.093750) ≈ 0.875000
			9'b001000100: sigmoid_out <= 9'b000011101;    //sigmoid(2.125000) ≈ 0.906250
			9'b001000101: sigmoid_out <= 9'b000011101;    //sigmoid(2.156250) ≈ 0.906250
			9'b001000110: sigmoid_out <= 9'b000011101;    //sigmoid(2.187500) ≈ 0.906250
			9'b001000111: sigmoid_out <= 9'b000011101;    //sigmoid(2.218750) ≈ 0.906250
			9'b001001000: sigmoid_out <= 9'b000011101;    //sigmoid(2.250000) ≈ 0.906250
			9'b001001001: sigmoid_out <= 9'b000011101;    //sigmoid(2.281250) ≈ 0.906250
			9'b001001010: sigmoid_out <= 9'b000011101;    //sigmoid(2.312500) ≈ 0.906250
			9'b001001011: sigmoid_out <= 9'b000011101;    //sigmoid(2.343750) ≈ 0.906250
			9'b001001100: sigmoid_out <= 9'b000011101;    //sigmoid(2.375000) ≈ 0.906250
			9'b001001101: sigmoid_out <= 9'b000011101;    //sigmoid(2.406250) ≈ 0.906250
			9'b001001110: sigmoid_out <= 9'b000011101;    //sigmoid(2.437500) ≈ 0.906250
			9'b001001111: sigmoid_out <= 9'b000011110;    //sigmoid(2.468750) ≈ 0.937500
			9'b001010000: sigmoid_out <= 9'b000011110;    //sigmoid(2.500000) ≈ 0.937500
			9'b001010001: sigmoid_out <= 9'b000011110;    //sigmoid(2.531250) ≈ 0.937500
			9'b001010010: sigmoid_out <= 9'b000011110;    //sigmoid(2.562500) ≈ 0.937500
			9'b001010011: sigmoid_out <= 9'b000011110;    //sigmoid(2.593750) ≈ 0.937500
			9'b001010100: sigmoid_out <= 9'b000011110;    //sigmoid(2.625000) ≈ 0.937500
			9'b001010101: sigmoid_out <= 9'b000011110;    //sigmoid(2.656250) ≈ 0.937500
			9'b001010110: sigmoid_out <= 9'b000011110;    //sigmoid(2.687500) ≈ 0.937500
			9'b001010111: sigmoid_out <= 9'b000011110;    //sigmoid(2.718750) ≈ 0.937500
			9'b001011000: sigmoid_out <= 9'b000011110;    //sigmoid(2.750000) ≈ 0.937500
			9'b001011001: sigmoid_out <= 9'b000011110;    //sigmoid(2.781250) ≈ 0.937500
			9'b001011010: sigmoid_out <= 9'b000011110;    //sigmoid(2.812500) ≈ 0.937500
			9'b001011011: sigmoid_out <= 9'b000011110;    //sigmoid(2.843750) ≈ 0.937500
			9'b001011100: sigmoid_out <= 9'b000011110;    //sigmoid(2.875000) ≈ 0.937500
			9'b001011101: sigmoid_out <= 9'b000011110;    //sigmoid(2.906250) ≈ 0.937500
			9'b001011110: sigmoid_out <= 9'b000011110;    //sigmoid(2.937500) ≈ 0.937500
			9'b001011111: sigmoid_out <= 9'b000011110;    //sigmoid(2.968750) ≈ 0.937500
			9'b001100000: sigmoid_out <= 9'b000011110;    //sigmoid(3.000000) ≈ 0.937500
			9'b001100001: sigmoid_out <= 9'b000011111;    //sigmoid(3.031250) ≈ 0.968750
			9'b001100010: sigmoid_out <= 9'b000011111;    //sigmoid(3.062500) ≈ 0.968750
			9'b001100011: sigmoid_out <= 9'b000011111;    //sigmoid(3.093750) ≈ 0.968750
			9'b001100100: sigmoid_out <= 9'b000011111;    //sigmoid(3.125000) ≈ 0.968750
			9'b001100101: sigmoid_out <= 9'b000011111;    //sigmoid(3.156250) ≈ 0.968750
			9'b001100110: sigmoid_out <= 9'b000011111;    //sigmoid(3.187500) ≈ 0.968750
			9'b001100111: sigmoid_out <= 9'b000011111;    //sigmoid(3.218750) ≈ 0.968750
			9'b001101000: sigmoid_out <= 9'b000011111;    //sigmoid(3.250000) ≈ 0.968750
			9'b001101001: sigmoid_out <= 9'b000011111;    //sigmoid(3.281250) ≈ 0.968750
			9'b001101010: sigmoid_out <= 9'b000011111;    //sigmoid(3.312500) ≈ 0.968750
			9'b001101011: sigmoid_out <= 9'b000011111;    //sigmoid(3.343750) ≈ 0.968750
			9'b001101100: sigmoid_out <= 9'b000011111;    //sigmoid(3.375000) ≈ 0.968750
			9'b001101101: sigmoid_out <= 9'b000011111;    //sigmoid(3.406250) ≈ 0.968750
			9'b001101110: sigmoid_out <= 9'b000011111;    //sigmoid(3.437500) ≈ 0.968750
			9'b001101111: sigmoid_out <= 9'b000011111;    //sigmoid(3.468750) ≈ 0.968750
			9'b001110000: sigmoid_out <= 9'b000011111;    //sigmoid(3.500000) ≈ 0.968750
			9'b001110001: sigmoid_out <= 9'b000011111;    //sigmoid(3.531250) ≈ 0.968750
			9'b001110010: sigmoid_out <= 9'b000011111;    //sigmoid(3.562500) ≈ 0.968750
			9'b001110011: sigmoid_out <= 9'b000011111;    //sigmoid(3.593750) ≈ 0.968750
			9'b001110100: sigmoid_out <= 9'b000011111;    //sigmoid(3.625000) ≈ 0.968750
			9'b001110101: sigmoid_out <= 9'b000011111;    //sigmoid(3.656250) ≈ 0.968750
			9'b001110110: sigmoid_out <= 9'b000011111;    //sigmoid(3.687500) ≈ 0.968750
			9'b001110111: sigmoid_out <= 9'b000011111;    //sigmoid(3.718750) ≈ 0.968750
			9'b001111000: sigmoid_out <= 9'b000011111;    //sigmoid(3.750000) ≈ 0.968750
			9'b001111001: sigmoid_out <= 9'b000011111;    //sigmoid(3.781250) ≈ 0.968750
			9'b001111010: sigmoid_out <= 9'b000011111;    //sigmoid(3.812500) ≈ 0.968750
			9'b001111011: sigmoid_out <= 9'b000011111;    //sigmoid(3.843750) ≈ 0.968750
			9'b001111100: sigmoid_out <= 9'b000011111;    //sigmoid(3.875000) ≈ 0.968750
			9'b001111101: sigmoid_out <= 9'b000011111;    //sigmoid(3.906250) ≈ 0.968750
			9'b001111110: sigmoid_out <= 9'b000011111;    //sigmoid(3.937500) ≈ 0.968750
			9'b001111111: sigmoid_out <= 9'b000011111;    //sigmoid(3.968750) ≈ 0.968750
			9'b010000000: sigmoid_out <= 9'b000011111;    //sigmoid(4.000000) ≈ 0.968750
			9'b010000001: sigmoid_out <= 9'b000011111;    //sigmoid(4.031250) ≈ 0.968750
			9'b010000010: sigmoid_out <= 9'b000011111;    //sigmoid(4.062500) ≈ 0.968750
			9'b010000011: sigmoid_out <= 9'b000011111;    //sigmoid(4.093750) ≈ 0.968750
			9'b010000100: sigmoid_out <= 9'b000011111;    //sigmoid(4.125000) ≈ 0.968750
			9'b010000101: sigmoid_out <= 9'b000100000;    //sigmoid(4.156250) ≈ 1.000000
			9'b010000110: sigmoid_out <= 9'b000100000;    //sigmoid(4.187500) ≈ 1.000000
			9'b010000111: sigmoid_out <= 9'b000100000;    //sigmoid(4.218750) ≈ 1.000000
			9'b010001000: sigmoid_out <= 9'b000100000;    //sigmoid(4.250000) ≈ 1.000000
			9'b010001001: sigmoid_out <= 9'b000100000;    //sigmoid(4.281250) ≈ 1.000000
			9'b010001010: sigmoid_out <= 9'b000100000;    //sigmoid(4.312500) ≈ 1.000000
			9'b010001011: sigmoid_out <= 9'b000100000;    //sigmoid(4.343750) ≈ 1.000000
			9'b010001100: sigmoid_out <= 9'b000100000;    //sigmoid(4.375000) ≈ 1.000000
			9'b010001101: sigmoid_out <= 9'b000100000;    //sigmoid(4.406250) ≈ 1.000000
			9'b010001110: sigmoid_out <= 9'b000100000;    //sigmoid(4.437500) ≈ 1.000000
			9'b010001111: sigmoid_out <= 9'b000100000;    //sigmoid(4.468750) ≈ 1.000000
			9'b010010000: sigmoid_out <= 9'b000100000;    //sigmoid(4.500000) ≈ 1.000000
			9'b010010001: sigmoid_out <= 9'b000100000;    //sigmoid(4.531250) ≈ 1.000000
			9'b010010010: sigmoid_out <= 9'b000100000;    //sigmoid(4.562500) ≈ 1.000000
			9'b010010011: sigmoid_out <= 9'b000100000;    //sigmoid(4.593750) ≈ 1.000000
			9'b010010100: sigmoid_out <= 9'b000100000;    //sigmoid(4.625000) ≈ 1.000000
			9'b010010101: sigmoid_out <= 9'b000100000;    //sigmoid(4.656250) ≈ 1.000000
			9'b010010110: sigmoid_out <= 9'b000100000;    //sigmoid(4.687500) ≈ 1.000000
			9'b010010111: sigmoid_out <= 9'b000100000;    //sigmoid(4.718750) ≈ 1.000000
			9'b010011000: sigmoid_out <= 9'b000100000;    //sigmoid(4.750000) ≈ 1.000000
			9'b010011001: sigmoid_out <= 9'b000100000;    //sigmoid(4.781250) ≈ 1.000000
			9'b010011010: sigmoid_out <= 9'b000100000;    //sigmoid(4.812500) ≈ 1.000000
			9'b010011011: sigmoid_out <= 9'b000100000;    //sigmoid(4.843750) ≈ 1.000000
			9'b010011100: sigmoid_out <= 9'b000100000;    //sigmoid(4.875000) ≈ 1.000000
			9'b010011101: sigmoid_out <= 9'b000100000;    //sigmoid(4.906250) ≈ 1.000000
			9'b010011110: sigmoid_out <= 9'b000100000;    //sigmoid(4.937500) ≈ 1.000000
			9'b010011111: sigmoid_out <= 9'b000100000;    //sigmoid(4.968750) ≈ 1.000000
			9'b010100000: sigmoid_out <= 9'b000100000;    //sigmoid(5.000000) ≈ 1.000000
			9'b010100001: sigmoid_out <= 9'b000100000;    //sigmoid(5.031250) ≈ 1.000000
			9'b010100010: sigmoid_out <= 9'b000100000;    //sigmoid(5.062500) ≈ 1.000000
			9'b010100011: sigmoid_out <= 9'b000100000;    //sigmoid(5.093750) ≈ 1.000000
			9'b010100100: sigmoid_out <= 9'b000100000;    //sigmoid(5.125000) ≈ 1.000000
			9'b010100101: sigmoid_out <= 9'b000100000;    //sigmoid(5.156250) ≈ 1.000000
			9'b010100110: sigmoid_out <= 9'b000100000;    //sigmoid(5.187500) ≈ 1.000000
			9'b010100111: sigmoid_out <= 9'b000100000;    //sigmoid(5.218750) ≈ 1.000000
			9'b010101000: sigmoid_out <= 9'b000100000;    //sigmoid(5.250000) ≈ 1.000000
			9'b010101001: sigmoid_out <= 9'b000100000;    //sigmoid(5.281250) ≈ 1.000000
			9'b010101010: sigmoid_out <= 9'b000100000;    //sigmoid(5.312500) ≈ 1.000000
			9'b010101011: sigmoid_out <= 9'b000100000;    //sigmoid(5.343750) ≈ 1.000000
			9'b010101100: sigmoid_out <= 9'b000100000;    //sigmoid(5.375000) ≈ 1.000000
			9'b010101101: sigmoid_out <= 9'b000100000;    //sigmoid(5.406250) ≈ 1.000000
			9'b010101110: sigmoid_out <= 9'b000100000;    //sigmoid(5.437500) ≈ 1.000000
			9'b010101111: sigmoid_out <= 9'b000100000;    //sigmoid(5.468750) ≈ 1.000000
			9'b010110000: sigmoid_out <= 9'b000100000;    //sigmoid(5.500000) ≈ 1.000000
			9'b010110001: sigmoid_out <= 9'b000100000;    //sigmoid(5.531250) ≈ 1.000000
			9'b010110010: sigmoid_out <= 9'b000100000;    //sigmoid(5.562500) ≈ 1.000000
			9'b010110011: sigmoid_out <= 9'b000100000;    //sigmoid(5.593750) ≈ 1.000000
			9'b010110100: sigmoid_out <= 9'b000100000;    //sigmoid(5.625000) ≈ 1.000000
			9'b010110101: sigmoid_out <= 9'b000100000;    //sigmoid(5.656250) ≈ 1.000000
			9'b010110110: sigmoid_out <= 9'b000100000;    //sigmoid(5.687500) ≈ 1.000000
			9'b010110111: sigmoid_out <= 9'b000100000;    //sigmoid(5.718750) ≈ 1.000000
			9'b010111000: sigmoid_out <= 9'b000100000;    //sigmoid(5.750000) ≈ 1.000000
			9'b010111001: sigmoid_out <= 9'b000100000;    //sigmoid(5.781250) ≈ 1.000000
			9'b010111010: sigmoid_out <= 9'b000100000;    //sigmoid(5.812500) ≈ 1.000000
			9'b010111011: sigmoid_out <= 9'b000100000;    //sigmoid(5.843750) ≈ 1.000000
			9'b010111100: sigmoid_out <= 9'b000100000;    //sigmoid(5.875000) ≈ 1.000000
			9'b010111101: sigmoid_out <= 9'b000100000;    //sigmoid(5.906250) ≈ 1.000000
			9'b010111110: sigmoid_out <= 9'b000100000;    //sigmoid(5.937500) ≈ 1.000000
			9'b010111111: sigmoid_out <= 9'b000100000;    //sigmoid(5.968750) ≈ 1.000000
			9'b011000000: sigmoid_out <= 9'b000100000;    //sigmoid(6.000000) ≈ 1.000000
			9'b011000001: sigmoid_out <= 9'b000100000;    //sigmoid(6.031250) ≈ 1.000000
			9'b011000010: sigmoid_out <= 9'b000100000;    //sigmoid(6.062500) ≈ 1.000000
			9'b011000011: sigmoid_out <= 9'b000100000;    //sigmoid(6.093750) ≈ 1.000000
			9'b011000100: sigmoid_out <= 9'b000100000;    //sigmoid(6.125000) ≈ 1.000000
			9'b011000101: sigmoid_out <= 9'b000100000;    //sigmoid(6.156250) ≈ 1.000000
			9'b011000110: sigmoid_out <= 9'b000100000;    //sigmoid(6.187500) ≈ 1.000000
			9'b011000111: sigmoid_out <= 9'b000100000;    //sigmoid(6.218750) ≈ 1.000000
			9'b011001000: sigmoid_out <= 9'b000100000;    //sigmoid(6.250000) ≈ 1.000000
			9'b011001001: sigmoid_out <= 9'b000100000;    //sigmoid(6.281250) ≈ 1.000000
			9'b011001010: sigmoid_out <= 9'b000100000;    //sigmoid(6.312500) ≈ 1.000000
			9'b011001011: sigmoid_out <= 9'b000100000;    //sigmoid(6.343750) ≈ 1.000000
			9'b011001100: sigmoid_out <= 9'b000100000;    //sigmoid(6.375000) ≈ 1.000000
			9'b011001101: sigmoid_out <= 9'b000100000;    //sigmoid(6.406250) ≈ 1.000000
			9'b011001110: sigmoid_out <= 9'b000100000;    //sigmoid(6.437500) ≈ 1.000000
			9'b011001111: sigmoid_out <= 9'b000100000;    //sigmoid(6.468750) ≈ 1.000000
			9'b011010000: sigmoid_out <= 9'b000100000;    //sigmoid(6.500000) ≈ 1.000000
			9'b011010001: sigmoid_out <= 9'b000100000;    //sigmoid(6.531250) ≈ 1.000000
			9'b011010010: sigmoid_out <= 9'b000100000;    //sigmoid(6.562500) ≈ 1.000000
			9'b011010011: sigmoid_out <= 9'b000100000;    //sigmoid(6.593750) ≈ 1.000000
			9'b011010100: sigmoid_out <= 9'b000100000;    //sigmoid(6.625000) ≈ 1.000000
			9'b011010101: sigmoid_out <= 9'b000100000;    //sigmoid(6.656250) ≈ 1.000000
			9'b011010110: sigmoid_out <= 9'b000100000;    //sigmoid(6.687500) ≈ 1.000000
			9'b011010111: sigmoid_out <= 9'b000100000;    //sigmoid(6.718750) ≈ 1.000000
			9'b011011000: sigmoid_out <= 9'b000100000;    //sigmoid(6.750000) ≈ 1.000000
			9'b011011001: sigmoid_out <= 9'b000100000;    //sigmoid(6.781250) ≈ 1.000000
			9'b011011010: sigmoid_out <= 9'b000100000;    //sigmoid(6.812500) ≈ 1.000000
			9'b011011011: sigmoid_out <= 9'b000100000;    //sigmoid(6.843750) ≈ 1.000000
			9'b011011100: sigmoid_out <= 9'b000100000;    //sigmoid(6.875000) ≈ 1.000000
			9'b011011101: sigmoid_out <= 9'b000100000;    //sigmoid(6.906250) ≈ 1.000000
			9'b011011110: sigmoid_out <= 9'b000100000;    //sigmoid(6.937500) ≈ 1.000000
			9'b011011111: sigmoid_out <= 9'b000100000;    //sigmoid(6.968750) ≈ 1.000000
			9'b011100000: sigmoid_out <= 9'b000100000;    //sigmoid(7.000000) ≈ 1.000000
			9'b011100001: sigmoid_out <= 9'b000100000;    //sigmoid(7.031250) ≈ 1.000000
			9'b011100010: sigmoid_out <= 9'b000100000;    //sigmoid(7.062500) ≈ 1.000000
			9'b011100011: sigmoid_out <= 9'b000100000;    //sigmoid(7.093750) ≈ 1.000000
			9'b011100100: sigmoid_out <= 9'b000100000;    //sigmoid(7.125000) ≈ 1.000000
			9'b011100101: sigmoid_out <= 9'b000100000;    //sigmoid(7.156250) ≈ 1.000000
			9'b011100110: sigmoid_out <= 9'b000100000;    //sigmoid(7.187500) ≈ 1.000000
			9'b011100111: sigmoid_out <= 9'b000100000;    //sigmoid(7.218750) ≈ 1.000000
			9'b011101000: sigmoid_out <= 9'b000100000;    //sigmoid(7.250000) ≈ 1.000000
			9'b011101001: sigmoid_out <= 9'b000100000;    //sigmoid(7.281250) ≈ 1.000000
			9'b011101010: sigmoid_out <= 9'b000100000;    //sigmoid(7.312500) ≈ 1.000000
			9'b011101011: sigmoid_out <= 9'b000100000;    //sigmoid(7.343750) ≈ 1.000000
			9'b011101100: sigmoid_out <= 9'b000100000;    //sigmoid(7.375000) ≈ 1.000000
			9'b011101101: sigmoid_out <= 9'b000100000;    //sigmoid(7.406250) ≈ 1.000000
			9'b011101110: sigmoid_out <= 9'b000100000;    //sigmoid(7.437500) ≈ 1.000000
			9'b011101111: sigmoid_out <= 9'b000100000;    //sigmoid(7.468750) ≈ 1.000000
			9'b011110000: sigmoid_out <= 9'b000100000;    //sigmoid(7.500000) ≈ 1.000000
			9'b011110001: sigmoid_out <= 9'b000100000;    //sigmoid(7.531250) ≈ 1.000000
			9'b011110010: sigmoid_out <= 9'b000100000;    //sigmoid(7.562500) ≈ 1.000000
			9'b011110011: sigmoid_out <= 9'b000100000;    //sigmoid(7.593750) ≈ 1.000000
			9'b011110100: sigmoid_out <= 9'b000100000;    //sigmoid(7.625000) ≈ 1.000000
			9'b011110101: sigmoid_out <= 9'b000100000;    //sigmoid(7.656250) ≈ 1.000000
			9'b011110110: sigmoid_out <= 9'b000100000;    //sigmoid(7.687500) ≈ 1.000000
			9'b011110111: sigmoid_out <= 9'b000100000;    //sigmoid(7.718750) ≈ 1.000000
			9'b011111000: sigmoid_out <= 9'b000100000;    //sigmoid(7.750000) ≈ 1.000000
			9'b011111001: sigmoid_out <= 9'b000100000;    //sigmoid(7.781250) ≈ 1.000000
			9'b011111010: sigmoid_out <= 9'b000100000;    //sigmoid(7.812500) ≈ 1.000000
			9'b011111011: sigmoid_out <= 9'b000100000;    //sigmoid(7.843750) ≈ 1.000000
			9'b011111100: sigmoid_out <= 9'b000100000;    //sigmoid(7.875000) ≈ 1.000000
			9'b011111101: sigmoid_out <= 9'b000100000;    //sigmoid(7.906250) ≈ 1.000000
			9'b011111110: sigmoid_out <= 9'b000100000;    //sigmoid(7.937500) ≈ 1.000000
			9'b011111111: sigmoid_out <= 9'b000100000;    //sigmoid(7.968750) ≈ 1.000000
			9'b100000000: sigmoid_out <= 9'b000100000;    //sigmoid(8.000000) ≈ 1.000000
			9'b100000001: sigmoid_out <= 9'b000100000;    //sigmoid(8.031250) ≈ 1.000000
			9'b100000010: sigmoid_out <= 9'b000100000;    //sigmoid(8.062500) ≈ 1.000000
			9'b100000011: sigmoid_out <= 9'b000100000;    //sigmoid(8.093750) ≈ 1.000000
			9'b100000100: sigmoid_out <= 9'b000100000;    //sigmoid(8.125000) ≈ 1.000000
			9'b100000101: sigmoid_out <= 9'b000100000;    //sigmoid(8.156250) ≈ 1.000000
			9'b100000110: sigmoid_out <= 9'b000100000;    //sigmoid(8.187500) ≈ 1.000000
			9'b100000111: sigmoid_out <= 9'b000100000;    //sigmoid(8.218750) ≈ 1.000000
			9'b100001000: sigmoid_out <= 9'b000100000;    //sigmoid(8.250000) ≈ 1.000000
			9'b100001001: sigmoid_out <= 9'b000100000;    //sigmoid(8.281250) ≈ 1.000000
			9'b100001010: sigmoid_out <= 9'b000100000;    //sigmoid(8.312500) ≈ 1.000000
			9'b100001011: sigmoid_out <= 9'b000100000;    //sigmoid(8.343750) ≈ 1.000000
			9'b100001100: sigmoid_out <= 9'b000100000;    //sigmoid(8.375000) ≈ 1.000000
			9'b100001101: sigmoid_out <= 9'b000100000;    //sigmoid(8.406250) ≈ 1.000000
			9'b100001110: sigmoid_out <= 9'b000100000;    //sigmoid(8.437500) ≈ 1.000000
			9'b100001111: sigmoid_out <= 9'b000100000;    //sigmoid(8.468750) ≈ 1.000000
			9'b100010000: sigmoid_out <= 9'b000100000;    //sigmoid(8.500000) ≈ 1.000000
			9'b100010001: sigmoid_out <= 9'b000100000;    //sigmoid(8.531250) ≈ 1.000000
			9'b100010010: sigmoid_out <= 9'b000100000;    //sigmoid(8.562500) ≈ 1.000000
			9'b100010011: sigmoid_out <= 9'b000100000;    //sigmoid(8.593750) ≈ 1.000000
			9'b100010100: sigmoid_out <= 9'b000100000;    //sigmoid(8.625000) ≈ 1.000000
			9'b100010101: sigmoid_out <= 9'b000100000;    //sigmoid(8.656250) ≈ 1.000000
			9'b100010110: sigmoid_out <= 9'b000100000;    //sigmoid(8.687500) ≈ 1.000000
			9'b100010111: sigmoid_out <= 9'b000100000;    //sigmoid(8.718750) ≈ 1.000000
			9'b100011000: sigmoid_out <= 9'b000100000;    //sigmoid(8.750000) ≈ 1.000000
			9'b100011001: sigmoid_out <= 9'b000100000;    //sigmoid(8.781250) ≈ 1.000000
			9'b100011010: sigmoid_out <= 9'b000100000;    //sigmoid(8.812500) ≈ 1.000000
			9'b100011011: sigmoid_out <= 9'b000100000;    //sigmoid(8.843750) ≈ 1.000000
			9'b100011100: sigmoid_out <= 9'b000100000;    //sigmoid(8.875000) ≈ 1.000000
			9'b100011101: sigmoid_out <= 9'b000100000;    //sigmoid(8.906250) ≈ 1.000000
			9'b100011110: sigmoid_out <= 9'b000100000;    //sigmoid(8.937500) ≈ 1.000000
			9'b100011111: sigmoid_out <= 9'b000100000;    //sigmoid(8.968750) ≈ 1.000000
			9'b100100000: sigmoid_out <= 9'b000100000;    //sigmoid(9.000000) ≈ 1.000000
			9'b100100001: sigmoid_out <= 9'b000100000;    //sigmoid(9.031250) ≈ 1.000000
			9'b100100010: sigmoid_out <= 9'b000100000;    //sigmoid(9.062500) ≈ 1.000000
			9'b100100011: sigmoid_out <= 9'b000100000;    //sigmoid(9.093750) ≈ 1.000000
			9'b100100100: sigmoid_out <= 9'b000100000;    //sigmoid(9.125000) ≈ 1.000000
			9'b100100101: sigmoid_out <= 9'b000100000;    //sigmoid(9.156250) ≈ 1.000000
			9'b100100110: sigmoid_out <= 9'b000100000;    //sigmoid(9.187500) ≈ 1.000000
			9'b100100111: sigmoid_out <= 9'b000100000;    //sigmoid(9.218750) ≈ 1.000000
			9'b100101000: sigmoid_out <= 9'b000100000;    //sigmoid(9.250000) ≈ 1.000000
			9'b100101001: sigmoid_out <= 9'b000100000;    //sigmoid(9.281250) ≈ 1.000000
			9'b100101010: sigmoid_out <= 9'b000100000;    //sigmoid(9.312500) ≈ 1.000000
			9'b100101011: sigmoid_out <= 9'b000100000;    //sigmoid(9.343750) ≈ 1.000000
			9'b100101100: sigmoid_out <= 9'b000100000;    //sigmoid(9.375000) ≈ 1.000000
			9'b100101101: sigmoid_out <= 9'b000100000;    //sigmoid(9.406250) ≈ 1.000000
			9'b100101110: sigmoid_out <= 9'b000100000;    //sigmoid(9.437500) ≈ 1.000000
			9'b100101111: sigmoid_out <= 9'b000100000;    //sigmoid(9.468750) ≈ 1.000000
			9'b100110000: sigmoid_out <= 9'b000100000;    //sigmoid(9.500000) ≈ 1.000000
			9'b100110001: sigmoid_out <= 9'b000100000;    //sigmoid(9.531250) ≈ 1.000000
			9'b100110010: sigmoid_out <= 9'b000100000;    //sigmoid(9.562500) ≈ 1.000000
			9'b100110011: sigmoid_out <= 9'b000100000;    //sigmoid(9.593750) ≈ 1.000000
			9'b100110100: sigmoid_out <= 9'b000100000;    //sigmoid(9.625000) ≈ 1.000000
			9'b100110101: sigmoid_out <= 9'b000100000;    //sigmoid(9.656250) ≈ 1.000000
			9'b100110110: sigmoid_out <= 9'b000100000;    //sigmoid(9.687500) ≈ 1.000000
			9'b100110111: sigmoid_out <= 9'b000100000;    //sigmoid(9.718750) ≈ 1.000000
			9'b100111000: sigmoid_out <= 9'b000100000;    //sigmoid(9.750000) ≈ 1.000000
			9'b100111001: sigmoid_out <= 9'b000100000;    //sigmoid(9.781250) ≈ 1.000000
			9'b100111010: sigmoid_out <= 9'b000100000;    //sigmoid(9.812500) ≈ 1.000000
			9'b100111011: sigmoid_out <= 9'b000100000;    //sigmoid(9.843750) ≈ 1.000000
			9'b100111100: sigmoid_out <= 9'b000100000;    //sigmoid(9.875000) ≈ 1.000000
			9'b100111101: sigmoid_out <= 9'b000100000;    //sigmoid(9.906250) ≈ 1.000000
			9'b100111110: sigmoid_out <= 9'b000100000;    //sigmoid(9.937500) ≈ 1.000000
			9'b100111111: sigmoid_out <= 9'b000100000;    //sigmoid(9.968750) ≈ 1.000000
			9'b101000000: sigmoid_out <= 9'b000100000;    //sigmoid(10.000000) ≈ 1.000000
			9'b101000001: sigmoid_out <= 9'b000100000;    //sigmoid(10.031250) ≈ 1.000000
			9'b101000010: sigmoid_out <= 9'b000100000;    //sigmoid(10.062500) ≈ 1.000000
			9'b101000011: sigmoid_out <= 9'b000100000;    //sigmoid(10.093750) ≈ 1.000000
			9'b101000100: sigmoid_out <= 9'b000100000;    //sigmoid(10.125000) ≈ 1.000000
			9'b101000101: sigmoid_out <= 9'b000100000;    //sigmoid(10.156250) ≈ 1.000000
			9'b101000110: sigmoid_out <= 9'b000100000;    //sigmoid(10.187500) ≈ 1.000000
			9'b101000111: sigmoid_out <= 9'b000100000;    //sigmoid(10.218750) ≈ 1.000000
			9'b101001000: sigmoid_out <= 9'b000100000;    //sigmoid(10.250000) ≈ 1.000000
			9'b101001001: sigmoid_out <= 9'b000100000;    //sigmoid(10.281250) ≈ 1.000000
			9'b101001010: sigmoid_out <= 9'b000100000;    //sigmoid(10.312500) ≈ 1.000000
			9'b101001011: sigmoid_out <= 9'b000100000;    //sigmoid(10.343750) ≈ 1.000000
			9'b101001100: sigmoid_out <= 9'b000100000;    //sigmoid(10.375000) ≈ 1.000000
			9'b101001101: sigmoid_out <= 9'b000100000;    //sigmoid(10.406250) ≈ 1.000000
			9'b101001110: sigmoid_out <= 9'b000100000;    //sigmoid(10.437500) ≈ 1.000000
			9'b101001111: sigmoid_out <= 9'b000100000;    //sigmoid(10.468750) ≈ 1.000000
			9'b101010000: sigmoid_out <= 9'b000100000;    //sigmoid(10.500000) ≈ 1.000000
			9'b101010001: sigmoid_out <= 9'b000100000;    //sigmoid(10.531250) ≈ 1.000000
			9'b101010010: sigmoid_out <= 9'b000100000;    //sigmoid(10.562500) ≈ 1.000000
			9'b101010011: sigmoid_out <= 9'b000100000;    //sigmoid(10.593750) ≈ 1.000000
			9'b101010100: sigmoid_out <= 9'b000100000;    //sigmoid(10.625000) ≈ 1.000000
			9'b101010101: sigmoid_out <= 9'b000100000;    //sigmoid(10.656250) ≈ 1.000000
			9'b101010110: sigmoid_out <= 9'b000100000;    //sigmoid(10.687500) ≈ 1.000000
			9'b101010111: sigmoid_out <= 9'b000100000;    //sigmoid(10.718750) ≈ 1.000000
			9'b101011000: sigmoid_out <= 9'b000100000;    //sigmoid(10.750000) ≈ 1.000000
			9'b101011001: sigmoid_out <= 9'b000100000;    //sigmoid(10.781250) ≈ 1.000000
			9'b101011010: sigmoid_out <= 9'b000100000;    //sigmoid(10.812500) ≈ 1.000000
			9'b101011011: sigmoid_out <= 9'b000100000;    //sigmoid(10.843750) ≈ 1.000000
			9'b101011100: sigmoid_out <= 9'b000100000;    //sigmoid(10.875000) ≈ 1.000000
			9'b101011101: sigmoid_out <= 9'b000100000;    //sigmoid(10.906250) ≈ 1.000000
			9'b101011110: sigmoid_out <= 9'b000100000;    //sigmoid(10.937500) ≈ 1.000000
			9'b101011111: sigmoid_out <= 9'b000100000;    //sigmoid(10.968750) ≈ 1.000000
			9'b101100000: sigmoid_out <= 9'b000100000;    //sigmoid(11.000000) ≈ 1.000000
			9'b101100001: sigmoid_out <= 9'b000100000;    //sigmoid(11.031250) ≈ 1.000000
			9'b101100010: sigmoid_out <= 9'b000100000;    //sigmoid(11.062500) ≈ 1.000000
			9'b101100011: sigmoid_out <= 9'b000100000;    //sigmoid(11.093750) ≈ 1.000000
			9'b101100100: sigmoid_out <= 9'b000100000;    //sigmoid(11.125000) ≈ 1.000000
			9'b101100101: sigmoid_out <= 9'b000100000;    //sigmoid(11.156250) ≈ 1.000000
			9'b101100110: sigmoid_out <= 9'b000100000;    //sigmoid(11.187500) ≈ 1.000000
			9'b101100111: sigmoid_out <= 9'b000100000;    //sigmoid(11.218750) ≈ 1.000000
			9'b101101000: sigmoid_out <= 9'b000100000;    //sigmoid(11.250000) ≈ 1.000000
			9'b101101001: sigmoid_out <= 9'b000100000;    //sigmoid(11.281250) ≈ 1.000000
			9'b101101010: sigmoid_out <= 9'b000100000;    //sigmoid(11.312500) ≈ 1.000000
			9'b101101011: sigmoid_out <= 9'b000100000;    //sigmoid(11.343750) ≈ 1.000000
			9'b101101100: sigmoid_out <= 9'b000100000;    //sigmoid(11.375000) ≈ 1.000000
			9'b101101101: sigmoid_out <= 9'b000100000;    //sigmoid(11.406250) ≈ 1.000000
			9'b101101110: sigmoid_out <= 9'b000100000;    //sigmoid(11.437500) ≈ 1.000000
			9'b101101111: sigmoid_out <= 9'b000100000;    //sigmoid(11.468750) ≈ 1.000000
			9'b101110000: sigmoid_out <= 9'b000100000;    //sigmoid(11.500000) ≈ 1.000000
			9'b101110001: sigmoid_out <= 9'b000100000;    //sigmoid(11.531250) ≈ 1.000000
			9'b101110010: sigmoid_out <= 9'b000100000;    //sigmoid(11.562500) ≈ 1.000000
			9'b101110011: sigmoid_out <= 9'b000100000;    //sigmoid(11.593750) ≈ 1.000000
			9'b101110100: sigmoid_out <= 9'b000100000;    //sigmoid(11.625000) ≈ 1.000000
			9'b101110101: sigmoid_out <= 9'b000100000;    //sigmoid(11.656250) ≈ 1.000000
			9'b101110110: sigmoid_out <= 9'b000100000;    //sigmoid(11.687500) ≈ 1.000000
			9'b101110111: sigmoid_out <= 9'b000100000;    //sigmoid(11.718750) ≈ 1.000000
			9'b101111000: sigmoid_out <= 9'b000100000;    //sigmoid(11.750000) ≈ 1.000000
			9'b101111001: sigmoid_out <= 9'b000100000;    //sigmoid(11.781250) ≈ 1.000000
			9'b101111010: sigmoid_out <= 9'b000100000;    //sigmoid(11.812500) ≈ 1.000000
			9'b101111011: sigmoid_out <= 9'b000100000;    //sigmoid(11.843750) ≈ 1.000000
			9'b101111100: sigmoid_out <= 9'b000100000;    //sigmoid(11.875000) ≈ 1.000000
			9'b101111101: sigmoid_out <= 9'b000100000;    //sigmoid(11.906250) ≈ 1.000000
			9'b101111110: sigmoid_out <= 9'b000100000;    //sigmoid(11.937500) ≈ 1.000000
			9'b101111111: sigmoid_out <= 9'b000100000;    //sigmoid(11.968750) ≈ 1.000000
			9'b110000000: sigmoid_out <= 9'b000100000;    //sigmoid(12.000000) ≈ 1.000000
			9'b110000001: sigmoid_out <= 9'b000100000;    //sigmoid(12.031250) ≈ 1.000000
			9'b110000010: sigmoid_out <= 9'b000100000;    //sigmoid(12.062500) ≈ 1.000000
			9'b110000011: sigmoid_out <= 9'b000100000;    //sigmoid(12.093750) ≈ 1.000000
			9'b110000100: sigmoid_out <= 9'b000100000;    //sigmoid(12.125000) ≈ 1.000000
			9'b110000101: sigmoid_out <= 9'b000100000;    //sigmoid(12.156250) ≈ 1.000000
			9'b110000110: sigmoid_out <= 9'b000100000;    //sigmoid(12.187500) ≈ 1.000000
			9'b110000111: sigmoid_out <= 9'b000100000;    //sigmoid(12.218750) ≈ 1.000000
			9'b110001000: sigmoid_out <= 9'b000100000;    //sigmoid(12.250000) ≈ 1.000000
			9'b110001001: sigmoid_out <= 9'b000100000;    //sigmoid(12.281250) ≈ 1.000000
			9'b110001010: sigmoid_out <= 9'b000100000;    //sigmoid(12.312500) ≈ 1.000000
			9'b110001011: sigmoid_out <= 9'b000100000;    //sigmoid(12.343750) ≈ 1.000000
			9'b110001100: sigmoid_out <= 9'b000100000;    //sigmoid(12.375000) ≈ 1.000000
			9'b110001101: sigmoid_out <= 9'b000100000;    //sigmoid(12.406250) ≈ 1.000000
			9'b110001110: sigmoid_out <= 9'b000100000;    //sigmoid(12.437500) ≈ 1.000000
			9'b110001111: sigmoid_out <= 9'b000100000;    //sigmoid(12.468750) ≈ 1.000000
			9'b110010000: sigmoid_out <= 9'b000100000;    //sigmoid(12.500000) ≈ 1.000000
			9'b110010001: sigmoid_out <= 9'b000100000;    //sigmoid(12.531250) ≈ 1.000000
			9'b110010010: sigmoid_out <= 9'b000100000;    //sigmoid(12.562500) ≈ 1.000000
			9'b110010011: sigmoid_out <= 9'b000100000;    //sigmoid(12.593750) ≈ 1.000000
			9'b110010100: sigmoid_out <= 9'b000100000;    //sigmoid(12.625000) ≈ 1.000000
			9'b110010101: sigmoid_out <= 9'b000100000;    //sigmoid(12.656250) ≈ 1.000000
			9'b110010110: sigmoid_out <= 9'b000100000;    //sigmoid(12.687500) ≈ 1.000000
			9'b110010111: sigmoid_out <= 9'b000100000;    //sigmoid(12.718750) ≈ 1.000000
			9'b110011000: sigmoid_out <= 9'b000100000;    //sigmoid(12.750000) ≈ 1.000000
			9'b110011001: sigmoid_out <= 9'b000100000;    //sigmoid(12.781250) ≈ 1.000000
			9'b110011010: sigmoid_out <= 9'b000100000;    //sigmoid(12.812500) ≈ 1.000000
			9'b110011011: sigmoid_out <= 9'b000100000;    //sigmoid(12.843750) ≈ 1.000000
			9'b110011100: sigmoid_out <= 9'b000100000;    //sigmoid(12.875000) ≈ 1.000000
			9'b110011101: sigmoid_out <= 9'b000100000;    //sigmoid(12.906250) ≈ 1.000000
			9'b110011110: sigmoid_out <= 9'b000100000;    //sigmoid(12.937500) ≈ 1.000000
			9'b110011111: sigmoid_out <= 9'b000100000;    //sigmoid(12.968750) ≈ 1.000000
			9'b110100000: sigmoid_out <= 9'b000100000;    //sigmoid(13.000000) ≈ 1.000000
			9'b110100001: sigmoid_out <= 9'b000100000;    //sigmoid(13.031250) ≈ 1.000000
			9'b110100010: sigmoid_out <= 9'b000100000;    //sigmoid(13.062500) ≈ 1.000000
			9'b110100011: sigmoid_out <= 9'b000100000;    //sigmoid(13.093750) ≈ 1.000000
			9'b110100100: sigmoid_out <= 9'b000100000;    //sigmoid(13.125000) ≈ 1.000000
			9'b110100101: sigmoid_out <= 9'b000100000;    //sigmoid(13.156250) ≈ 1.000000
			9'b110100110: sigmoid_out <= 9'b000100000;    //sigmoid(13.187500) ≈ 1.000000
			9'b110100111: sigmoid_out <= 9'b000100000;    //sigmoid(13.218750) ≈ 1.000000
			9'b110101000: sigmoid_out <= 9'b000100000;    //sigmoid(13.250000) ≈ 1.000000
			9'b110101001: sigmoid_out <= 9'b000100000;    //sigmoid(13.281250) ≈ 1.000000
			9'b110101010: sigmoid_out <= 9'b000100000;    //sigmoid(13.312500) ≈ 1.000000
			9'b110101011: sigmoid_out <= 9'b000100000;    //sigmoid(13.343750) ≈ 1.000000
			9'b110101100: sigmoid_out <= 9'b000100000;    //sigmoid(13.375000) ≈ 1.000000
			9'b110101101: sigmoid_out <= 9'b000100000;    //sigmoid(13.406250) ≈ 1.000000
			9'b110101110: sigmoid_out <= 9'b000100000;    //sigmoid(13.437500) ≈ 1.000000
			9'b110101111: sigmoid_out <= 9'b000100000;    //sigmoid(13.468750) ≈ 1.000000
			9'b110110000: sigmoid_out <= 9'b000100000;    //sigmoid(13.500000) ≈ 1.000000
			9'b110110001: sigmoid_out <= 9'b000100000;    //sigmoid(13.531250) ≈ 1.000000
			9'b110110010: sigmoid_out <= 9'b000100000;    //sigmoid(13.562500) ≈ 1.000000
			9'b110110011: sigmoid_out <= 9'b000100000;    //sigmoid(13.593750) ≈ 1.000000
			9'b110110100: sigmoid_out <= 9'b000100000;    //sigmoid(13.625000) ≈ 1.000000
			9'b110110101: sigmoid_out <= 9'b000100000;    //sigmoid(13.656250) ≈ 1.000000
			9'b110110110: sigmoid_out <= 9'b000100000;    //sigmoid(13.687500) ≈ 1.000000
			9'b110110111: sigmoid_out <= 9'b000100000;    //sigmoid(13.718750) ≈ 1.000000
			9'b110111000: sigmoid_out <= 9'b000100000;    //sigmoid(13.750000) ≈ 1.000000
			9'b110111001: sigmoid_out <= 9'b000100000;    //sigmoid(13.781250) ≈ 1.000000
			9'b110111010: sigmoid_out <= 9'b000100000;    //sigmoid(13.812500) ≈ 1.000000
			9'b110111011: sigmoid_out <= 9'b000100000;    //sigmoid(13.843750) ≈ 1.000000
			9'b110111100: sigmoid_out <= 9'b000100000;    //sigmoid(13.875000) ≈ 1.000000
			9'b110111101: sigmoid_out <= 9'b000100000;    //sigmoid(13.906250) ≈ 1.000000
			9'b110111110: sigmoid_out <= 9'b000100000;    //sigmoid(13.937500) ≈ 1.000000
			9'b110111111: sigmoid_out <= 9'b000100000;    //sigmoid(13.968750) ≈ 1.000000
			9'b111000000: sigmoid_out <= 9'b000100000;    //sigmoid(14.000000) ≈ 1.000000
			9'b111000001: sigmoid_out <= 9'b000100000;    //sigmoid(14.031250) ≈ 1.000000
			9'b111000010: sigmoid_out <= 9'b000100000;    //sigmoid(14.062500) ≈ 1.000000
			9'b111000011: sigmoid_out <= 9'b000100000;    //sigmoid(14.093750) ≈ 1.000000
			9'b111000100: sigmoid_out <= 9'b000100000;    //sigmoid(14.125000) ≈ 1.000000
			9'b111000101: sigmoid_out <= 9'b000100000;    //sigmoid(14.156250) ≈ 1.000000
			9'b111000110: sigmoid_out <= 9'b000100000;    //sigmoid(14.187500) ≈ 1.000000
			9'b111000111: sigmoid_out <= 9'b000100000;    //sigmoid(14.218750) ≈ 1.000000
			9'b111001000: sigmoid_out <= 9'b000100000;    //sigmoid(14.250000) ≈ 1.000000
			9'b111001001: sigmoid_out <= 9'b000100000;    //sigmoid(14.281250) ≈ 1.000000
			9'b111001010: sigmoid_out <= 9'b000100000;    //sigmoid(14.312500) ≈ 1.000000
			9'b111001011: sigmoid_out <= 9'b000100000;    //sigmoid(14.343750) ≈ 1.000000
			9'b111001100: sigmoid_out <= 9'b000100000;    //sigmoid(14.375000) ≈ 1.000000
			9'b111001101: sigmoid_out <= 9'b000100000;    //sigmoid(14.406250) ≈ 1.000000
			9'b111001110: sigmoid_out <= 9'b000100000;    //sigmoid(14.437500) ≈ 1.000000
			9'b111001111: sigmoid_out <= 9'b000100000;    //sigmoid(14.468750) ≈ 1.000000
			9'b111010000: sigmoid_out <= 9'b000100000;    //sigmoid(14.500000) ≈ 1.000000
			9'b111010001: sigmoid_out <= 9'b000100000;    //sigmoid(14.531250) ≈ 1.000000
			9'b111010010: sigmoid_out <= 9'b000100000;    //sigmoid(14.562500) ≈ 1.000000
			9'b111010011: sigmoid_out <= 9'b000100000;    //sigmoid(14.593750) ≈ 1.000000
			9'b111010100: sigmoid_out <= 9'b000100000;    //sigmoid(14.625000) ≈ 1.000000
			9'b111010101: sigmoid_out <= 9'b000100000;    //sigmoid(14.656250) ≈ 1.000000
			9'b111010110: sigmoid_out <= 9'b000100000;    //sigmoid(14.687500) ≈ 1.000000
			9'b111010111: sigmoid_out <= 9'b000100000;    //sigmoid(14.718750) ≈ 1.000000
			9'b111011000: sigmoid_out <= 9'b000100000;    //sigmoid(14.750000) ≈ 1.000000
			9'b111011001: sigmoid_out <= 9'b000100000;    //sigmoid(14.781250) ≈ 1.000000
			9'b111011010: sigmoid_out <= 9'b000100000;    //sigmoid(14.812500) ≈ 1.000000
			9'b111011011: sigmoid_out <= 9'b000100000;    //sigmoid(14.843750) ≈ 1.000000
			9'b111011100: sigmoid_out <= 9'b000100000;    //sigmoid(14.875000) ≈ 1.000000
			9'b111011101: sigmoid_out <= 9'b000100000;    //sigmoid(14.906250) ≈ 1.000000
			9'b111011110: sigmoid_out <= 9'b000100000;    //sigmoid(14.937500) ≈ 1.000000
			9'b111011111: sigmoid_out <= 9'b000100000;    //sigmoid(14.968750) ≈ 1.000000
			9'b111100000: sigmoid_out <= 9'b000100000;    //sigmoid(15.000000) ≈ 1.000000
			9'b111100001: sigmoid_out <= 9'b000100000;    //sigmoid(15.031250) ≈ 1.000000
			9'b111100010: sigmoid_out <= 9'b000100000;    //sigmoid(15.062500) ≈ 1.000000
			9'b111100011: sigmoid_out <= 9'b000100000;    //sigmoid(15.093750) ≈ 1.000000
			9'b111100100: sigmoid_out <= 9'b000100000;    //sigmoid(15.125000) ≈ 1.000000
			9'b111100101: sigmoid_out <= 9'b000100000;    //sigmoid(15.156250) ≈ 1.000000
			9'b111100110: sigmoid_out <= 9'b000100000;    //sigmoid(15.187500) ≈ 1.000000
			9'b111100111: sigmoid_out <= 9'b000100000;    //sigmoid(15.218750) ≈ 1.000000
			9'b111101000: sigmoid_out <= 9'b000100000;    //sigmoid(15.250000) ≈ 1.000000
			9'b111101001: sigmoid_out <= 9'b000100000;    //sigmoid(15.281250) ≈ 1.000000
			9'b111101010: sigmoid_out <= 9'b000100000;    //sigmoid(15.312500) ≈ 1.000000
			9'b111101011: sigmoid_out <= 9'b000100000;    //sigmoid(15.343750) ≈ 1.000000
			9'b111101100: sigmoid_out <= 9'b000100000;    //sigmoid(15.375000) ≈ 1.000000
			9'b111101101: sigmoid_out <= 9'b000100000;    //sigmoid(15.406250) ≈ 1.000000
			9'b111101110: sigmoid_out <= 9'b000100000;    //sigmoid(15.437500) ≈ 1.000000
			9'b111101111: sigmoid_out <= 9'b000100000;    //sigmoid(15.468750) ≈ 1.000000
			9'b111110000: sigmoid_out <= 9'b000100000;    //sigmoid(15.500000) ≈ 1.000000
			9'b111110001: sigmoid_out <= 9'b000100000;    //sigmoid(15.531250) ≈ 1.000000
			9'b111110010: sigmoid_out <= 9'b000100000;    //sigmoid(15.562500) ≈ 1.000000
			9'b111110011: sigmoid_out <= 9'b000100000;    //sigmoid(15.593750) ≈ 1.000000
			9'b111110100: sigmoid_out <= 9'b000100000;    //sigmoid(15.625000) ≈ 1.000000
			9'b111110101: sigmoid_out <= 9'b000100000;    //sigmoid(15.656250) ≈ 1.000000
			9'b111110110: sigmoid_out <= 9'b000100000;    //sigmoid(15.687500) ≈ 1.000000
			9'b111110111: sigmoid_out <= 9'b000100000;    //sigmoid(15.718750) ≈ 1.000000
			9'b111111000: sigmoid_out <= 9'b000100000;    //sigmoid(15.750000) ≈ 1.000000
			9'b111111001: sigmoid_out <= 9'b000100000;    //sigmoid(15.781250) ≈ 1.000000
			9'b111111010: sigmoid_out <= 9'b000100000;    //sigmoid(15.812500) ≈ 1.000000
			9'b111111011: sigmoid_out <= 9'b000100000;    //sigmoid(15.843750) ≈ 1.000000
			9'b111111100: sigmoid_out <= 9'b000100000;    //sigmoid(15.875000) ≈ 1.000000
			9'b111111101: sigmoid_out <= 9'b000100000;    //sigmoid(15.906250) ≈ 1.000000
			9'b111111110: sigmoid_out <= 9'b000100000;    //sigmoid(15.937500) ≈ 1.000000
			9'b111111111: sigmoid_out <= 9'b000100000;    //sigmoid(15.968750) ≈ 1.000000

        endcase
    end
endmodule