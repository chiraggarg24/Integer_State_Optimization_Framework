//////////////////////////////////////////////////////////////////////////////////
// Company: LEED
// Engineer: Philip Canoza
// 
// Create Date: 2019-06-28 12:04:12.135005
// Design Name: vanilla
// Module Name: sigmoidLUT_8bit_6point
// Project Name: RBM_FPGA
// Description: An implementation of a sigmoid function via 8 bit LUT.
//              It is assumed that all inputs are unsigned fixed point values.
// 
// Additional Comments: Generated by LUT_generator_sigmoid.py
// 
//////////////////////////////////////////////////////////////////////////////////
module sigmoidLUT_8bit_6point #(
    parameter PRECISION_BITS = 8
)(
    input[PRECISION_BITS - 1: 0] sigmoid_in,
    output reg[PRECISION_BITS - 1: 0] sigmoid_out
);

    always @(sigmoid_in) begin
        case(sigmoid_in)
			8'b00000000: sigmoid_out <= 8'b00100000;    //sigmoid(0.000000) ≈ 0.500000
			8'b00000001: sigmoid_out <= 8'b00100000;    //sigmoid(0.015625) ≈ 0.500000
			8'b00000010: sigmoid_out <= 8'b00100000;    //sigmoid(0.031250) ≈ 0.500000
			8'b00000011: sigmoid_out <= 8'b00100001;    //sigmoid(0.046875) ≈ 0.515625
			8'b00000100: sigmoid_out <= 8'b00100001;    //sigmoid(0.062500) ≈ 0.515625
			8'b00000101: sigmoid_out <= 8'b00100001;    //sigmoid(0.078125) ≈ 0.515625
			8'b00000110: sigmoid_out <= 8'b00100001;    //sigmoid(0.093750) ≈ 0.515625
			8'b00000111: sigmoid_out <= 8'b00100010;    //sigmoid(0.109375) ≈ 0.531250
			8'b00001000: sigmoid_out <= 8'b00100010;    //sigmoid(0.125000) ≈ 0.531250
			8'b00001001: sigmoid_out <= 8'b00100010;    //sigmoid(0.140625) ≈ 0.531250
			8'b00001010: sigmoid_out <= 8'b00100010;    //sigmoid(0.156250) ≈ 0.531250
			8'b00001011: sigmoid_out <= 8'b00100011;    //sigmoid(0.171875) ≈ 0.546875
			8'b00001100: sigmoid_out <= 8'b00100011;    //sigmoid(0.187500) ≈ 0.546875
			8'b00001101: sigmoid_out <= 8'b00100011;    //sigmoid(0.203125) ≈ 0.546875
			8'b00001110: sigmoid_out <= 8'b00100011;    //sigmoid(0.218750) ≈ 0.546875
			8'b00001111: sigmoid_out <= 8'b00100100;    //sigmoid(0.234375) ≈ 0.562500
			8'b00010000: sigmoid_out <= 8'b00100100;    //sigmoid(0.250000) ≈ 0.562500
			8'b00010001: sigmoid_out <= 8'b00100100;    //sigmoid(0.265625) ≈ 0.562500
			8'b00010010: sigmoid_out <= 8'b00100100;    //sigmoid(0.281250) ≈ 0.562500
			8'b00010011: sigmoid_out <= 8'b00100101;    //sigmoid(0.296875) ≈ 0.578125
			8'b00010100: sigmoid_out <= 8'b00100101;    //sigmoid(0.312500) ≈ 0.578125
			8'b00010101: sigmoid_out <= 8'b00100101;    //sigmoid(0.328125) ≈ 0.578125
			8'b00010110: sigmoid_out <= 8'b00100101;    //sigmoid(0.343750) ≈ 0.578125
			8'b00010111: sigmoid_out <= 8'b00100110;    //sigmoid(0.359375) ≈ 0.593750
			8'b00011000: sigmoid_out <= 8'b00100110;    //sigmoid(0.375000) ≈ 0.593750
			8'b00011001: sigmoid_out <= 8'b00100110;    //sigmoid(0.390625) ≈ 0.593750
			8'b00011010: sigmoid_out <= 8'b00100110;    //sigmoid(0.406250) ≈ 0.593750
			8'b00011011: sigmoid_out <= 8'b00100111;    //sigmoid(0.421875) ≈ 0.609375
			8'b00011100: sigmoid_out <= 8'b00100111;    //sigmoid(0.437500) ≈ 0.609375
			8'b00011101: sigmoid_out <= 8'b00100111;    //sigmoid(0.453125) ≈ 0.609375
			8'b00011110: sigmoid_out <= 8'b00100111;    //sigmoid(0.468750) ≈ 0.609375
			8'b00011111: sigmoid_out <= 8'b00101000;    //sigmoid(0.484375) ≈ 0.625000
			8'b00100000: sigmoid_out <= 8'b00101000;    //sigmoid(0.500000) ≈ 0.625000
			8'b00100001: sigmoid_out <= 8'b00101000;    //sigmoid(0.515625) ≈ 0.625000
			8'b00100010: sigmoid_out <= 8'b00101000;    //sigmoid(0.531250) ≈ 0.625000
			8'b00100011: sigmoid_out <= 8'b00101001;    //sigmoid(0.546875) ≈ 0.640625
			8'b00100100: sigmoid_out <= 8'b00101001;    //sigmoid(0.562500) ≈ 0.640625
			8'b00100101: sigmoid_out <= 8'b00101001;    //sigmoid(0.578125) ≈ 0.640625
			8'b00100110: sigmoid_out <= 8'b00101001;    //sigmoid(0.593750) ≈ 0.640625
			8'b00100111: sigmoid_out <= 8'b00101001;    //sigmoid(0.609375) ≈ 0.640625
			8'b00101000: sigmoid_out <= 8'b00101010;    //sigmoid(0.625000) ≈ 0.656250
			8'b00101001: sigmoid_out <= 8'b00101010;    //sigmoid(0.640625) ≈ 0.656250
			8'b00101010: sigmoid_out <= 8'b00101010;    //sigmoid(0.656250) ≈ 0.656250
			8'b00101011: sigmoid_out <= 8'b00101010;    //sigmoid(0.671875) ≈ 0.656250
			8'b00101100: sigmoid_out <= 8'b00101011;    //sigmoid(0.687500) ≈ 0.671875
			8'b00101101: sigmoid_out <= 8'b00101011;    //sigmoid(0.703125) ≈ 0.671875
			8'b00101110: sigmoid_out <= 8'b00101011;    //sigmoid(0.718750) ≈ 0.671875
			8'b00101111: sigmoid_out <= 8'b00101011;    //sigmoid(0.734375) ≈ 0.671875
			8'b00110000: sigmoid_out <= 8'b00101011;    //sigmoid(0.750000) ≈ 0.671875
			8'b00110001: sigmoid_out <= 8'b00101100;    //sigmoid(0.765625) ≈ 0.687500
			8'b00110010: sigmoid_out <= 8'b00101100;    //sigmoid(0.781250) ≈ 0.687500
			8'b00110011: sigmoid_out <= 8'b00101100;    //sigmoid(0.796875) ≈ 0.687500
			8'b00110100: sigmoid_out <= 8'b00101100;    //sigmoid(0.812500) ≈ 0.687500
			8'b00110101: sigmoid_out <= 8'b00101101;    //sigmoid(0.828125) ≈ 0.703125
			8'b00110110: sigmoid_out <= 8'b00101101;    //sigmoid(0.843750) ≈ 0.703125
			8'b00110111: sigmoid_out <= 8'b00101101;    //sigmoid(0.859375) ≈ 0.703125
			8'b00111000: sigmoid_out <= 8'b00101101;    //sigmoid(0.875000) ≈ 0.703125
			8'b00111001: sigmoid_out <= 8'b00101101;    //sigmoid(0.890625) ≈ 0.703125
			8'b00111010: sigmoid_out <= 8'b00101110;    //sigmoid(0.906250) ≈ 0.718750
			8'b00111011: sigmoid_out <= 8'b00101110;    //sigmoid(0.921875) ≈ 0.718750
			8'b00111100: sigmoid_out <= 8'b00101110;    //sigmoid(0.937500) ≈ 0.718750
			8'b00111101: sigmoid_out <= 8'b00101110;    //sigmoid(0.953125) ≈ 0.718750
			8'b00111110: sigmoid_out <= 8'b00101110;    //sigmoid(0.968750) ≈ 0.718750
			8'b00111111: sigmoid_out <= 8'b00101111;    //sigmoid(0.984375) ≈ 0.734375
			8'b01000000: sigmoid_out <= 8'b00101111;    //sigmoid(1.000000) ≈ 0.734375
			8'b01000001: sigmoid_out <= 8'b00101111;    //sigmoid(1.015625) ≈ 0.734375
			8'b01000010: sigmoid_out <= 8'b00101111;    //sigmoid(1.031250) ≈ 0.734375
			8'b01000011: sigmoid_out <= 8'b00101111;    //sigmoid(1.046875) ≈ 0.734375
			8'b01000100: sigmoid_out <= 8'b00110000;    //sigmoid(1.062500) ≈ 0.750000
			8'b01000101: sigmoid_out <= 8'b00110000;    //sigmoid(1.078125) ≈ 0.750000
			8'b01000110: sigmoid_out <= 8'b00110000;    //sigmoid(1.093750) ≈ 0.750000
			8'b01000111: sigmoid_out <= 8'b00110000;    //sigmoid(1.109375) ≈ 0.750000
			8'b01001000: sigmoid_out <= 8'b00110000;    //sigmoid(1.125000) ≈ 0.750000
			8'b01001001: sigmoid_out <= 8'b00110000;    //sigmoid(1.140625) ≈ 0.750000
			8'b01001010: sigmoid_out <= 8'b00110001;    //sigmoid(1.156250) ≈ 0.765625
			8'b01001011: sigmoid_out <= 8'b00110001;    //sigmoid(1.171875) ≈ 0.765625
			8'b01001100: sigmoid_out <= 8'b00110001;    //sigmoid(1.187500) ≈ 0.765625
			8'b01001101: sigmoid_out <= 8'b00110001;    //sigmoid(1.203125) ≈ 0.765625
			8'b01001110: sigmoid_out <= 8'b00110001;    //sigmoid(1.218750) ≈ 0.765625
			8'b01001111: sigmoid_out <= 8'b00110010;    //sigmoid(1.234375) ≈ 0.781250
			8'b01010000: sigmoid_out <= 8'b00110010;    //sigmoid(1.250000) ≈ 0.781250
			8'b01010001: sigmoid_out <= 8'b00110010;    //sigmoid(1.265625) ≈ 0.781250
			8'b01010010: sigmoid_out <= 8'b00110010;    //sigmoid(1.281250) ≈ 0.781250
			8'b01010011: sigmoid_out <= 8'b00110010;    //sigmoid(1.296875) ≈ 0.781250
			8'b01010100: sigmoid_out <= 8'b00110010;    //sigmoid(1.312500) ≈ 0.781250
			8'b01010101: sigmoid_out <= 8'b00110011;    //sigmoid(1.328125) ≈ 0.796875
			8'b01010110: sigmoid_out <= 8'b00110011;    //sigmoid(1.343750) ≈ 0.796875
			8'b01010111: sigmoid_out <= 8'b00110011;    //sigmoid(1.359375) ≈ 0.796875
			8'b01011000: sigmoid_out <= 8'b00110011;    //sigmoid(1.375000) ≈ 0.796875
			8'b01011001: sigmoid_out <= 8'b00110011;    //sigmoid(1.390625) ≈ 0.796875
			8'b01011010: sigmoid_out <= 8'b00110011;    //sigmoid(1.406250) ≈ 0.796875
			8'b01011011: sigmoid_out <= 8'b00110100;    //sigmoid(1.421875) ≈ 0.812500
			8'b01011100: sigmoid_out <= 8'b00110100;    //sigmoid(1.437500) ≈ 0.812500
			8'b01011101: sigmoid_out <= 8'b00110100;    //sigmoid(1.453125) ≈ 0.812500
			8'b01011110: sigmoid_out <= 8'b00110100;    //sigmoid(1.468750) ≈ 0.812500
			8'b01011111: sigmoid_out <= 8'b00110100;    //sigmoid(1.484375) ≈ 0.812500
			8'b01100000: sigmoid_out <= 8'b00110100;    //sigmoid(1.500000) ≈ 0.812500
			8'b01100001: sigmoid_out <= 8'b00110100;    //sigmoid(1.515625) ≈ 0.812500
			8'b01100010: sigmoid_out <= 8'b00110101;    //sigmoid(1.531250) ≈ 0.828125
			8'b01100011: sigmoid_out <= 8'b00110101;    //sigmoid(1.546875) ≈ 0.828125
			8'b01100100: sigmoid_out <= 8'b00110101;    //sigmoid(1.562500) ≈ 0.828125
			8'b01100101: sigmoid_out <= 8'b00110101;    //sigmoid(1.578125) ≈ 0.828125
			8'b01100110: sigmoid_out <= 8'b00110101;    //sigmoid(1.593750) ≈ 0.828125
			8'b01100111: sigmoid_out <= 8'b00110101;    //sigmoid(1.609375) ≈ 0.828125
			8'b01101000: sigmoid_out <= 8'b00110101;    //sigmoid(1.625000) ≈ 0.828125
			8'b01101001: sigmoid_out <= 8'b00110110;    //sigmoid(1.640625) ≈ 0.843750
			8'b01101010: sigmoid_out <= 8'b00110110;    //sigmoid(1.656250) ≈ 0.843750
			8'b01101011: sigmoid_out <= 8'b00110110;    //sigmoid(1.671875) ≈ 0.843750
			8'b01101100: sigmoid_out <= 8'b00110110;    //sigmoid(1.687500) ≈ 0.843750
			8'b01101101: sigmoid_out <= 8'b00110110;    //sigmoid(1.703125) ≈ 0.843750
			8'b01101110: sigmoid_out <= 8'b00110110;    //sigmoid(1.718750) ≈ 0.843750
			8'b01101111: sigmoid_out <= 8'b00110110;    //sigmoid(1.734375) ≈ 0.843750
			8'b01110000: sigmoid_out <= 8'b00110111;    //sigmoid(1.750000) ≈ 0.859375
			8'b01110001: sigmoid_out <= 8'b00110111;    //sigmoid(1.765625) ≈ 0.859375
			8'b01110010: sigmoid_out <= 8'b00110111;    //sigmoid(1.781250) ≈ 0.859375
			8'b01110011: sigmoid_out <= 8'b00110111;    //sigmoid(1.796875) ≈ 0.859375
			8'b01110100: sigmoid_out <= 8'b00110111;    //sigmoid(1.812500) ≈ 0.859375
			8'b01110101: sigmoid_out <= 8'b00110111;    //sigmoid(1.828125) ≈ 0.859375
			8'b01110110: sigmoid_out <= 8'b00110111;    //sigmoid(1.843750) ≈ 0.859375
			8'b01110111: sigmoid_out <= 8'b00110111;    //sigmoid(1.859375) ≈ 0.859375
			8'b01111000: sigmoid_out <= 8'b00110111;    //sigmoid(1.875000) ≈ 0.859375
			8'b01111001: sigmoid_out <= 8'b00111000;    //sigmoid(1.890625) ≈ 0.875000
			8'b01111010: sigmoid_out <= 8'b00111000;    //sigmoid(1.906250) ≈ 0.875000
			8'b01111011: sigmoid_out <= 8'b00111000;    //sigmoid(1.921875) ≈ 0.875000
			8'b01111100: sigmoid_out <= 8'b00111000;    //sigmoid(1.937500) ≈ 0.875000
			8'b01111101: sigmoid_out <= 8'b00111000;    //sigmoid(1.953125) ≈ 0.875000
			8'b01111110: sigmoid_out <= 8'b00111000;    //sigmoid(1.968750) ≈ 0.875000
			8'b01111111: sigmoid_out <= 8'b00111000;    //sigmoid(1.984375) ≈ 0.875000
			8'b10000000: sigmoid_out <= 8'b00111000;    //sigmoid(2.000000) ≈ 0.875000
			8'b10000001: sigmoid_out <= 8'b00111000;    //sigmoid(2.015625) ≈ 0.875000
			8'b10000010: sigmoid_out <= 8'b00111001;    //sigmoid(2.031250) ≈ 0.890625
			8'b10000011: sigmoid_out <= 8'b00111001;    //sigmoid(2.046875) ≈ 0.890625
			8'b10000100: sigmoid_out <= 8'b00111001;    //sigmoid(2.062500) ≈ 0.890625
			8'b10000101: sigmoid_out <= 8'b00111001;    //sigmoid(2.078125) ≈ 0.890625
			8'b10000110: sigmoid_out <= 8'b00111001;    //sigmoid(2.093750) ≈ 0.890625
			8'b10000111: sigmoid_out <= 8'b00111001;    //sigmoid(2.109375) ≈ 0.890625
			8'b10001000: sigmoid_out <= 8'b00111001;    //sigmoid(2.125000) ≈ 0.890625
			8'b10001001: sigmoid_out <= 8'b00111001;    //sigmoid(2.140625) ≈ 0.890625
			8'b10001010: sigmoid_out <= 8'b00111001;    //sigmoid(2.156250) ≈ 0.890625
			8'b10001011: sigmoid_out <= 8'b00111001;    //sigmoid(2.171875) ≈ 0.890625
			8'b10001100: sigmoid_out <= 8'b00111010;    //sigmoid(2.187500) ≈ 0.906250
			8'b10001101: sigmoid_out <= 8'b00111010;    //sigmoid(2.203125) ≈ 0.906250
			8'b10001110: sigmoid_out <= 8'b00111010;    //sigmoid(2.218750) ≈ 0.906250
			8'b10001111: sigmoid_out <= 8'b00111010;    //sigmoid(2.234375) ≈ 0.906250
			8'b10010000: sigmoid_out <= 8'b00111010;    //sigmoid(2.250000) ≈ 0.906250
			8'b10010001: sigmoid_out <= 8'b00111010;    //sigmoid(2.265625) ≈ 0.906250
			8'b10010010: sigmoid_out <= 8'b00111010;    //sigmoid(2.281250) ≈ 0.906250
			8'b10010011: sigmoid_out <= 8'b00111010;    //sigmoid(2.296875) ≈ 0.906250
			8'b10010100: sigmoid_out <= 8'b00111010;    //sigmoid(2.312500) ≈ 0.906250
			8'b10010101: sigmoid_out <= 8'b00111010;    //sigmoid(2.328125) ≈ 0.906250
			8'b10010110: sigmoid_out <= 8'b00111010;    //sigmoid(2.343750) ≈ 0.906250
			8'b10010111: sigmoid_out <= 8'b00111010;    //sigmoid(2.359375) ≈ 0.906250
			8'b10011000: sigmoid_out <= 8'b00111011;    //sigmoid(2.375000) ≈ 0.921875
			8'b10011001: sigmoid_out <= 8'b00111011;    //sigmoid(2.390625) ≈ 0.921875
			8'b10011010: sigmoid_out <= 8'b00111011;    //sigmoid(2.406250) ≈ 0.921875
			8'b10011011: sigmoid_out <= 8'b00111011;    //sigmoid(2.421875) ≈ 0.921875
			8'b10011100: sigmoid_out <= 8'b00111011;    //sigmoid(2.437500) ≈ 0.921875
			8'b10011101: sigmoid_out <= 8'b00111011;    //sigmoid(2.453125) ≈ 0.921875
			8'b10011110: sigmoid_out <= 8'b00111011;    //sigmoid(2.468750) ≈ 0.921875
			8'b10011111: sigmoid_out <= 8'b00111011;    //sigmoid(2.484375) ≈ 0.921875
			8'b10100000: sigmoid_out <= 8'b00111011;    //sigmoid(2.500000) ≈ 0.921875
			8'b10100001: sigmoid_out <= 8'b00111011;    //sigmoid(2.515625) ≈ 0.921875
			8'b10100010: sigmoid_out <= 8'b00111011;    //sigmoid(2.531250) ≈ 0.921875
			8'b10100011: sigmoid_out <= 8'b00111011;    //sigmoid(2.546875) ≈ 0.921875
			8'b10100100: sigmoid_out <= 8'b00111011;    //sigmoid(2.562500) ≈ 0.921875
			8'b10100101: sigmoid_out <= 8'b00111011;    //sigmoid(2.578125) ≈ 0.921875
			8'b10100110: sigmoid_out <= 8'b00111100;    //sigmoid(2.593750) ≈ 0.937500
			8'b10100111: sigmoid_out <= 8'b00111100;    //sigmoid(2.609375) ≈ 0.937500
			8'b10101000: sigmoid_out <= 8'b00111100;    //sigmoid(2.625000) ≈ 0.937500
			8'b10101001: sigmoid_out <= 8'b00111100;    //sigmoid(2.640625) ≈ 0.937500
			8'b10101010: sigmoid_out <= 8'b00111100;    //sigmoid(2.656250) ≈ 0.937500
			8'b10101011: sigmoid_out <= 8'b00111100;    //sigmoid(2.671875) ≈ 0.937500
			8'b10101100: sigmoid_out <= 8'b00111100;    //sigmoid(2.687500) ≈ 0.937500
			8'b10101101: sigmoid_out <= 8'b00111100;    //sigmoid(2.703125) ≈ 0.937500
			8'b10101110: sigmoid_out <= 8'b00111100;    //sigmoid(2.718750) ≈ 0.937500
			8'b10101111: sigmoid_out <= 8'b00111100;    //sigmoid(2.734375) ≈ 0.937500
			8'b10110000: sigmoid_out <= 8'b00111100;    //sigmoid(2.750000) ≈ 0.937500
			8'b10110001: sigmoid_out <= 8'b00111100;    //sigmoid(2.765625) ≈ 0.937500
			8'b10110010: sigmoid_out <= 8'b00111100;    //sigmoid(2.781250) ≈ 0.937500
			8'b10110011: sigmoid_out <= 8'b00111100;    //sigmoid(2.796875) ≈ 0.937500
			8'b10110100: sigmoid_out <= 8'b00111100;    //sigmoid(2.812500) ≈ 0.937500
			8'b10110101: sigmoid_out <= 8'b00111100;    //sigmoid(2.828125) ≈ 0.937500
			8'b10110110: sigmoid_out <= 8'b00111100;    //sigmoid(2.843750) ≈ 0.937500
			8'b10110111: sigmoid_out <= 8'b00111101;    //sigmoid(2.859375) ≈ 0.953125
			8'b10111000: sigmoid_out <= 8'b00111101;    //sigmoid(2.875000) ≈ 0.953125
			8'b10111001: sigmoid_out <= 8'b00111101;    //sigmoid(2.890625) ≈ 0.953125
			8'b10111010: sigmoid_out <= 8'b00111101;    //sigmoid(2.906250) ≈ 0.953125
			8'b10111011: sigmoid_out <= 8'b00111101;    //sigmoid(2.921875) ≈ 0.953125
			8'b10111100: sigmoid_out <= 8'b00111101;    //sigmoid(2.937500) ≈ 0.953125
			8'b10111101: sigmoid_out <= 8'b00111101;    //sigmoid(2.953125) ≈ 0.953125
			8'b10111110: sigmoid_out <= 8'b00111101;    //sigmoid(2.968750) ≈ 0.953125
			8'b10111111: sigmoid_out <= 8'b00111101;    //sigmoid(2.984375) ≈ 0.953125
			8'b11000000: sigmoid_out <= 8'b00111101;    //sigmoid(3.000000) ≈ 0.953125
			8'b11000001: sigmoid_out <= 8'b00111101;    //sigmoid(3.015625) ≈ 0.953125
			8'b11000010: sigmoid_out <= 8'b00111101;    //sigmoid(3.031250) ≈ 0.953125
			8'b11000011: sigmoid_out <= 8'b00111101;    //sigmoid(3.046875) ≈ 0.953125
			8'b11000100: sigmoid_out <= 8'b00111101;    //sigmoid(3.062500) ≈ 0.953125
			8'b11000101: sigmoid_out <= 8'b00111101;    //sigmoid(3.078125) ≈ 0.953125
			8'b11000110: sigmoid_out <= 8'b00111101;    //sigmoid(3.093750) ≈ 0.953125
			8'b11000111: sigmoid_out <= 8'b00111101;    //sigmoid(3.109375) ≈ 0.953125
			8'b11001000: sigmoid_out <= 8'b00111101;    //sigmoid(3.125000) ≈ 0.953125
			8'b11001001: sigmoid_out <= 8'b00111101;    //sigmoid(3.140625) ≈ 0.953125
			8'b11001010: sigmoid_out <= 8'b00111101;    //sigmoid(3.156250) ≈ 0.953125
			8'b11001011: sigmoid_out <= 8'b00111101;    //sigmoid(3.171875) ≈ 0.953125
			8'b11001100: sigmoid_out <= 8'b00111101;    //sigmoid(3.187500) ≈ 0.953125
			8'b11001101: sigmoid_out <= 8'b00111110;    //sigmoid(3.203125) ≈ 0.968750
			8'b11001110: sigmoid_out <= 8'b00111110;    //sigmoid(3.218750) ≈ 0.968750
			8'b11001111: sigmoid_out <= 8'b00111110;    //sigmoid(3.234375) ≈ 0.968750
			8'b11010000: sigmoid_out <= 8'b00111110;    //sigmoid(3.250000) ≈ 0.968750
			8'b11010001: sigmoid_out <= 8'b00111110;    //sigmoid(3.265625) ≈ 0.968750
			8'b11010010: sigmoid_out <= 8'b00111110;    //sigmoid(3.281250) ≈ 0.968750
			8'b11010011: sigmoid_out <= 8'b00111110;    //sigmoid(3.296875) ≈ 0.968750
			8'b11010100: sigmoid_out <= 8'b00111110;    //sigmoid(3.312500) ≈ 0.968750
			8'b11010101: sigmoid_out <= 8'b00111110;    //sigmoid(3.328125) ≈ 0.968750
			8'b11010110: sigmoid_out <= 8'b00111110;    //sigmoid(3.343750) ≈ 0.968750
			8'b11010111: sigmoid_out <= 8'b00111110;    //sigmoid(3.359375) ≈ 0.968750
			8'b11011000: sigmoid_out <= 8'b00111110;    //sigmoid(3.375000) ≈ 0.968750
			8'b11011001: sigmoid_out <= 8'b00111110;    //sigmoid(3.390625) ≈ 0.968750
			8'b11011010: sigmoid_out <= 8'b00111110;    //sigmoid(3.406250) ≈ 0.968750
			8'b11011011: sigmoid_out <= 8'b00111110;    //sigmoid(3.421875) ≈ 0.968750
			8'b11011100: sigmoid_out <= 8'b00111110;    //sigmoid(3.437500) ≈ 0.968750
			8'b11011101: sigmoid_out <= 8'b00111110;    //sigmoid(3.453125) ≈ 0.968750
			8'b11011110: sigmoid_out <= 8'b00111110;    //sigmoid(3.468750) ≈ 0.968750
			8'b11011111: sigmoid_out <= 8'b00111110;    //sigmoid(3.484375) ≈ 0.968750
			8'b11100000: sigmoid_out <= 8'b00111110;    //sigmoid(3.500000) ≈ 0.968750
			8'b11100001: sigmoid_out <= 8'b00111110;    //sigmoid(3.515625) ≈ 0.968750
			8'b11100010: sigmoid_out <= 8'b00111110;    //sigmoid(3.531250) ≈ 0.968750
			8'b11100011: sigmoid_out <= 8'b00111110;    //sigmoid(3.546875) ≈ 0.968750
			8'b11100100: sigmoid_out <= 8'b00111110;    //sigmoid(3.562500) ≈ 0.968750
			8'b11100101: sigmoid_out <= 8'b00111110;    //sigmoid(3.578125) ≈ 0.968750
			8'b11100110: sigmoid_out <= 8'b00111110;    //sigmoid(3.593750) ≈ 0.968750
			8'b11100111: sigmoid_out <= 8'b00111110;    //sigmoid(3.609375) ≈ 0.968750
			8'b11101000: sigmoid_out <= 8'b00111110;    //sigmoid(3.625000) ≈ 0.968750
			8'b11101001: sigmoid_out <= 8'b00111110;    //sigmoid(3.640625) ≈ 0.968750
			8'b11101010: sigmoid_out <= 8'b00111110;    //sigmoid(3.656250) ≈ 0.968750
			8'b11101011: sigmoid_out <= 8'b00111110;    //sigmoid(3.671875) ≈ 0.968750
			8'b11101100: sigmoid_out <= 8'b00111110;    //sigmoid(3.687500) ≈ 0.968750
			8'b11101101: sigmoid_out <= 8'b00111110;    //sigmoid(3.703125) ≈ 0.968750
			8'b11101110: sigmoid_out <= 8'b00111110;    //sigmoid(3.718750) ≈ 0.968750
			8'b11101111: sigmoid_out <= 8'b00111111;    //sigmoid(3.734375) ≈ 0.984375
			8'b11110000: sigmoid_out <= 8'b00111111;    //sigmoid(3.750000) ≈ 0.984375
			8'b11110001: sigmoid_out <= 8'b00111111;    //sigmoid(3.765625) ≈ 0.984375
			8'b11110010: sigmoid_out <= 8'b00111111;    //sigmoid(3.781250) ≈ 0.984375
			8'b11110011: sigmoid_out <= 8'b00111111;    //sigmoid(3.796875) ≈ 0.984375
			8'b11110100: sigmoid_out <= 8'b00111111;    //sigmoid(3.812500) ≈ 0.984375
			8'b11110101: sigmoid_out <= 8'b00111111;    //sigmoid(3.828125) ≈ 0.984375
			8'b11110110: sigmoid_out <= 8'b00111111;    //sigmoid(3.843750) ≈ 0.984375
			8'b11110111: sigmoid_out <= 8'b00111111;    //sigmoid(3.859375) ≈ 0.984375
			8'b11111000: sigmoid_out <= 8'b00111111;    //sigmoid(3.875000) ≈ 0.984375
			8'b11111001: sigmoid_out <= 8'b00111111;    //sigmoid(3.890625) ≈ 0.984375
			8'b11111010: sigmoid_out <= 8'b00111111;    //sigmoid(3.906250) ≈ 0.984375
			8'b11111011: sigmoid_out <= 8'b00111111;    //sigmoid(3.921875) ≈ 0.984375
			8'b11111100: sigmoid_out <= 8'b00111111;    //sigmoid(3.937500) ≈ 0.984375
			8'b11111101: sigmoid_out <= 8'b00111111;    //sigmoid(3.953125) ≈ 0.984375
			8'b11111110: sigmoid_out <= 8'b00111111;    //sigmoid(3.968750) ≈ 0.984375
			8'b11111111: sigmoid_out <= 8'b00111111;    //sigmoid(3.984375) ≈ 0.984375

        endcase
    end
endmodule